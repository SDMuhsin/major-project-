`timescale 1ns / 1ps
module Function_generator1 (f,adrs,rst);
parameter K_N=1022;
parameter addr_width=4;
output reg [K_N-1:0]f;
input [addr_width-1:0]adrs;
input rst;
input rst;
always@(adrs,rst)begin
  if(rst)begin
    f = K_N'd0;
  end
  else begin
    case(adrs)begin
    addr_width'd0 : begin 
      f = K_N'b10111010110011100101010110111111010101101100110001010101001010000011110111111110111011111110101010001100100011001111111100000100111000011110101111011001000001100111011100010000100110001000111000100101000001001000110101100111010100100101010000100110100100111001111000100000011010001101001011011100011011111100110100101111100000100010101111101011011010111101100101101100100010100111011011110100100100110010101010101110100110111100010100111010110100100000101000101010100111001000011010111011010001100001111001000010010111010010100011010000101010110101110000010000110100110001010010100001010101000110000010100010111011010000111100100111101110000100011100001010100010010101111001111111110100110000111001110010001000000100001101010101111011000111000001110100110010100000011010000001001110000111100111010010111000110101000000010110011111011001110000100100011011000111110111010000000100110100000000111011001000100100000010011110001100000010001000100100011111010101011100001100111110100111110010000001110100011000110010100100101100;
    end 
    addr_width'd1 : begin 
      f = K_N'b01100010101100100001110011110000101011101110000001100100100111111010011001111011011111010000111010100110010101010001110000011100110100011001010011001010011101110101000000011110000011111100111110001100100001011000011001111011100111001111011001111001110000011000101111001111011110010011100111100001000011111000010101010000011001100001100001001000101001001110000010101001111010011110110110110111110110101011100111101101101010111010000110001100000101101000110010001110001010001010101011001101110111101010101100011110110010010110111000111110100100001101010110101010111000100100101011001100000110001000101000100100010010001111011001000101001111100000000000101111011101001100100100111000110110000010001000101001000111110110000000010110111000010000000100000101000011011110001101010010111100100000111010010001101001010010110101001011001001111111010010011111101001011000110110101111010101011110111011101010000111100001100011100011011001100011010111011100101101101000000000011000111111101011101011100111010101011110000000001110001000;
    end 
    addr_width'd2 : begin 
      f = K_N'b01101000000110101000111001010001010000100000101111011000001010010100111011001110000100111110010010010001110101100001100000001000001111111111101110111010100000110000110110110101111110101111001100110000001000001001100001110111110110000000000111111001001010110101111000000111000100010111110001010111111001110101111101101111000011011000011100111011001111100101001000001111001000011110101011111101011110001100000101100001001011000110001000101000000100010001101000110110100111010101011110010000111101011001001010011010000010011011111000111011101011101111111000111000010000011000001111110110101011100001101011111011101011110100001001000011001111010101110110011101010010010110010100001110111001010000010011001010001101100001111111111100111000100111101111100110011100010100110001100100110001110111100000011100011001001001010100001111110001011011100000110101101011001001100100111110001000010101010101001011000010111101101011010010000010110010100011011101110000101100111101001110011110011110000010010101101001010101111100100100001100;
    end 
    addr_width'd3 : begin 
      f = K_N'b00110101100101010001111111101110011011110010000011001001000000100010100101101100100101001000100000000000001100110100010111100110110001010101001001101100010101010001100100100011000001000101010011000101010101101011100010100000010011111100000011011100011001000010110101101000001011011001010010110100010110010100101101010001100101110000001101111101111100010101101101011000000101111011001001101111000101101101000010100011001100000010110000001001001110000011010000010010100000100010111101101101001010110010001101001110111011010000001110011110111111100100111100000111000000011100010100011110001001001100010101100100010111101000000101111110011010000000101101111111011100100100011000100011010100010100011010011010000100001001100000010000110010001100100011101110111010000110001110110111111110111011101001011101000001010100010111001100111010000101011101011010110010100110011101101010001101100101011110111101110000000110111011111101001111101101110011000111101110010100000101100001111000111011111100101111110011100111101010111001101100;
    end 
    addr_width'd4 : begin 
      f = K_N'b00011000100000010101011110101110010000011000001100000111010001001011101011100000101011011010011000101001010111100000100010110111100110100100010000001000000111100001000100011111011010011011101111100111100000110001110100000111101111101110101111110111011000100011001011100000011001011111011101010010110101001111001000011000110100111001101101101100010110111111001000001010111001011011100011111111000101110010101001111111000111110110100000001110011010111111010110101010110000111100010000110100001101110011011011000010101110110000000101001100000000001111100000101110101101101011100000011011101100010001010010001000010010001000000111000101100001010011100011010100001001101101011101111001110000011011001010110100101100010101000001110110100100011001010000011100111010001110100111010010100011101101100100100101110001100111101000101100100101111111111100101000011101001100001110011100001000000110001110111111111010001000001101100001011000101110101001000001001101101001001100000111001010011110100011110010100011001000100001110010010111;
    end 
    addr_width'd5 : begin 
      f = K_N'b01100000110011010001111100011100001010000010101000010110000100100110010101111110100011000111110000010100001000000011001100101100101000100100010111000000011101010110111101111000011101000100110010000000011110010110011011000011111000010011001001100100001110001000011110001011110100101100110011001000001100111000100001000001010110100110000100100111000001011010101100011001001010110011010100010010111011101111000011011001010100100100100011110111101101110011111001011011000011110100000100101011111101110110110110110100100001101001011011010010111101110011000110010011111001111100100100001010000001011001000110110111101100010010001110100001010000000111000011010011001011000010100011011011110101111101111000100011101010010111000001100110000001100111110000001011110110111000010100011111000000010001111001001011110100011110011000101000001001101011110011001100111010110110111011000001000101101100110111101111111111100110011100100100011000010000010010000101001001100000000001001011101110111000100101110110110010111001101011110110110111;
    end 
    addr_width'd6 : begin 
      f = K_N'b01110110011010000101010100010010010111001111110111001000000001001101101011111000110110111110001101100110000011101000011010000110010000100000001000110000111011010100111000000100100111011111000100011101100000101110001101010111110001010100111111100010010101101110101000000001111101010110100000011101100101010101010001001100011110100001111000110010101101111100001100001010100011100110110011110101110100001000011010011110011101010100111111111101111001101010111011111010011011010111101111101000111100011011000101001000010001000101001011101011101001100100101101001001000011111111110010101100000101001101101000101000110001100010001010101111000110110011100010101010000000111010010100010111100000010100001111110110100100011001001101111011010000101110011111010000110100100010011001110100011101010101001010100000110110001000010101011101001111101000110011011101000010101100001000111111100010111111000111101110100111001000011100101100011100011010110011011010010111100000000110001101000001010011000011110101001011011011000100010000111110;
    end 
    addr_width'd7 : begin 
      f = K_N'b00010100101101011111100110001110100011010101010111111100100011101001101101001110111001000101001111000110100101100011111000000101001000010100011110101000010101111010110000011110000010000110011101011101100110011010001100001000111001110010011010011111101011000101011000000000110101111011000101010101110111101000110010110001101110101100011110000110111101000101101101000110101101010010001100000111001101101001001011011110011101000101111111011111000100000111001001001101110110100011100011111101000010010011101100011100001101101110001101011111111101110000001000101111011110011111000101101011101000000000010101010011001111111101110101001001001010100000011110000000011010110011011000001010110100101100011111111100101001001110001000101000000111001100010011011110110111110001111110011101001111100101001101100110111000001000111111110011100101010001001111010111100111001110110000001000000010111000110001001110111111100110010100100000110010111011111001000011010101100111011011101111001101010110011111010001100100010010101010101000000000;
    end 
    addr_width'd8 : begin 
      f = K_N'b00000000000010001011010011101000100110011110010111110111111001101001001010111101110011100110100111001110001111111010110110011001011100011000001111001111101011101011001001111000010111010000110000111101100111001010111001010001000000110001011011010100101111010110010110100010101000000110110010111010011111110100111001001100010010101000000010000011100110101100101010000001000000010010001101000011011001001000111011101010100011011011101110100010010001100100101001101000111000010001010110101011001111110100000000110100101101101111111111001101000000010001010000100001110101001000010111111101111000011101101100110110100000110010010000011111000001000000010001100001000010111000001000001101111101110111100000111110101011010110101011001111010000101000010010101110000001000011011110001011111110110100110000011001011101000000101101100001000111110101101011011011100001110110000010000010000001010010101100010000100110001111100110011011110000011100101011000110100011111010110010010011101111001101101110111001110111010110000110010010101111;
    end 
    addr_width'd9 : begin 
      f = K_N'b01011110100110110010101100110011111011111000001011010000111001100100101010100010001000100110110101101010000010101101110011010001011110011101010110010011001011101110000111001111010000000001101100110011011001000100100111010000111111110111011101010111010101001100101001010110011001010000011100010110111001100001101001000011111110010110001111010101100110000110010111000111111100000001011111110101001110000011000001010001010000110000011001100100100110000010001011001010101001110010110000010101001011110110111010110010010110011011000000101000000110010001010001101111101111000001101000000100110000100100101100111110110001110101010001010100100001000001010100011111000000111111110110010110110011000011101101110100101110001100010110111110110110010000001011110110100101001100001110100101011110000011111000001101000101001010000110111111101000011101010100011111110000110111101001110000111011000000001000001100010111000100010011101101010010010011000011110100001100110100111000010110100011000001100010101001111001000010101111000011000010;
    end 
    addr_width'd10 : begin 
      f = K_N'b00000110111100011111111100100100100100011001001011110010111010101111000001100011010010001000111000100110011111101110111010011001010011100111011101100000100110010101110001001111101001101111111110100000111001000010010000011000001001011010011111110101101101100101110001110100111110110001011010101100010011001000100100011011110000000000100011010011001110101101010011111111100101110101001000111110111001011011110100010100000100100110100100010110111000000101000000101111111100101111100011100100101000000111111111000010110010100101000011110000100000011010000000000100100001100100111100011110100000111001110000100010101011011010001100001101000111100100100111000000010111110010001110100111010000110001000011010101100111010010000011011001110011101000001011001100010101101000000101101001110111111011111101110010000111101110110110000011010110111011000100001001101100100100000101011111010100010110011010000100111111011101011100001001010011101011001111110100000001011100000000001100011010101110100001111110101000010111001010000101111000;
    end 
    addr_width'd11 : begin 
      f = K_N'b01000001000010011101101000101010001001001110010000011011000111110011011101010110010001010010001010011001100000011101010010110111111010001000110000110110101000010010110110101011011001001110100100011100011101100100110011000100001111001100111011000001100010001110110010001100010110000101010111001000111111110100100010001011101110010001000000000011011000000010101111101111010000111101101111101100010010100110001000010000010010001001000001101010001011001101110001011101101111010100000100000011010000110001110110111000010000110000101111000111011110001110000011101101011101001010001101010101101011010110001100110011100100011000110000010111100110101110000111010000010010001011011100001110100100100100111000100110110111001101101100011011101010100100111110111110000011010010011110111000001000010100001110010001110010100011011010110111110100100111111111101110101001110001111101000010011100010110011001101010111001110001111010000110001010100110110000110101011111110001100011100111011111101000000010110010011101011100010001010111110010;
    end 
    addr_width'd12 : begin 
      f = K_N'b00100010100010000100010101110111010110100010011000100101000001011011010001110010100010001110000001100101101100100011101101001010011011010111100010101111101111011101101100100011010101101011001110010010110001101001001011101111010101101010001101011010101101001010101000100111011101100111110111100111001011110000010110001100011001001000010001000101011111001001010110101000110011001101110100001110111100100010010110101011101001010110101101110110010101111011011111110000111010010100011111011100000101111111100101110010010011000110000110001101111011110011000011110001110010100001100111101011010101111010011010100111010011011101101100000001011111010101100110001110001011010010001011110011110101001010111010000110101111001000100010000010001101111000111110101010110011000010011011011011111101010011000001100000001100111110011010001000011110111101000111001001100011000001001010000001011110001001110001100011101110011101010110101010001010011010111010101011010111110010101101001100010001001011000010111010110100101010111001001101001001;
    end 
    addr_width'd13 : begin 
      f = K_N'b01110010011100111110100000110100001010010001100011100000100101111011000111000001111101011111111011110011001010100001010100001010111011110101111000010001000110000100011110000010101101011011110101011010000111011000000001110001111010010100010101111000101100001010110001110010001011010111101111110100100111101000110001111000110100111001000100101001010000110111000111111111101110100111101110001000111110101011111110001100110000000011101001100010101110010100000011001110011000001101011001101001110111111011011110110110000100001111110101000010010000001000010011110010011001100000111000001000101101100101000001111010111001100000101111010010011110110001111011101000111001001010000001101001110011101111101001001011101001111111111000001000011101011011100010111111000101101011011000110000110110110110111000010101001011010001010100000010110100000110101111011111011010101110101100101010010111010101110011111101010010011100111011011011111000011010101111100001001011101011001000011100001101000101010100101111000000000100101010101110011111;
    end 
default: f = K_N'd0;    endcase
  end
  endmodule
