`timescale 1ns / 1ps
module LMem1To0_511_circ13_combined_ys_yu_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        rxIn,
        load_input_en,
        iteration_0_indicator,
        feedback_en,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter r_lower = 32;
parameter c = 17;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input load_input_en;
input iteration_0_indicator;
input [ADDRESSWIDTH-1:0]unloadAddress;
input feedback_en;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input [ r_lower * w - 1 : 0 ] rxIn; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
wire [w-1:0]rxInConnector[r_lower-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

generate
    for (k=0;k<r_lower;k=k+1)begin:assign_rx
        assign rxInConnector[k] = rxIn[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            if(feedback_en)begin
                 fifoOut[i][0] <= fifoOut[i][c-1];
            end
            else if(load_input_en)begin
                 if(i < r_lower)begin
                   fifoOut[i][0] = rxInConnector[i];
                 end
                 else begin
                   fifoOut[i][0] = maxVal;
                 end
            end
            else begin
                 fifoOut[i][0] <= ly0InConnector[i];
            end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
       0: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = fifoOut[17][14][w-1];
              unloadMuxOut[20] = fifoOut[18][14][w-1];
              unloadMuxOut[21] = fifoOut[19][14][w-1];
              unloadMuxOut[22] = fifoOut[20][14][w-1];
              unloadMuxOut[23] = fifoOut[21][14][w-1];
              unloadMuxOut[24] = fifoOut[22][14][w-1];
              unloadMuxOut[25] = fifoOut[23][14][w-1];
              unloadMuxOut[26] = fifoOut[24][14][w-1];
              unloadMuxOut[27] = fifoOut[25][14][w-1];
              unloadMuxOut[28] = fifoOut[0][13][w-1];
              unloadMuxOut[29] = fifoOut[1][13][w-1];
              unloadMuxOut[30] = fifoOut[2][13][w-1];
              unloadMuxOut[31] = fifoOut[3][13][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[4][14][w-1];
              unloadMuxOut[1] = fifoOut[5][14][w-1];
              unloadMuxOut[2] = fifoOut[6][14][w-1];
              unloadMuxOut[3] = fifoOut[7][14][w-1];
              unloadMuxOut[4] = fifoOut[8][14][w-1];
              unloadMuxOut[5] = fifoOut[9][14][w-1];
              unloadMuxOut[6] = fifoOut[10][14][w-1];
              unloadMuxOut[7] = fifoOut[11][14][w-1];
              unloadMuxOut[8] = fifoOut[12][14][w-1];
              unloadMuxOut[9] = fifoOut[13][14][w-1];
              unloadMuxOut[10] = fifoOut[14][14][w-1];
              unloadMuxOut[11] = fifoOut[15][14][w-1];
              unloadMuxOut[12] = fifoOut[16][14][w-1];
              unloadMuxOut[13] = fifoOut[17][14][w-1];
              unloadMuxOut[14] = fifoOut[18][14][w-1];
              unloadMuxOut[15] = fifoOut[19][14][w-1];
              unloadMuxOut[16] = fifoOut[20][14][w-1];
              unloadMuxOut[17] = fifoOut[21][14][w-1];
              unloadMuxOut[18] = fifoOut[22][14][w-1];
              unloadMuxOut[19] = fifoOut[23][14][w-1];
              unloadMuxOut[20] = fifoOut[24][14][w-1];
              unloadMuxOut[21] = fifoOut[25][14][w-1];
              unloadMuxOut[22] = fifoOut[0][13][w-1];
              unloadMuxOut[23] = fifoOut[1][13][w-1];
              unloadMuxOut[24] = fifoOut[2][13][w-1];
              unloadMuxOut[25] = fifoOut[3][13][w-1];
              unloadMuxOut[26] = fifoOut[4][13][w-1];
              unloadMuxOut[27] = fifoOut[5][13][w-1];
              unloadMuxOut[28] = fifoOut[6][13][w-1];
              unloadMuxOut[29] = fifoOut[7][13][w-1];
              unloadMuxOut[30] = fifoOut[8][13][w-1];
              unloadMuxOut[31] = fifoOut[9][13][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[10][14][w-1];
              unloadMuxOut[1] = fifoOut[11][14][w-1];
              unloadMuxOut[2] = fifoOut[12][14][w-1];
              unloadMuxOut[3] = fifoOut[13][14][w-1];
              unloadMuxOut[4] = fifoOut[14][14][w-1];
              unloadMuxOut[5] = fifoOut[15][14][w-1];
              unloadMuxOut[6] = fifoOut[16][14][w-1];
              unloadMuxOut[7] = fifoOut[17][14][w-1];
              unloadMuxOut[8] = fifoOut[18][14][w-1];
              unloadMuxOut[9] = fifoOut[19][14][w-1];
              unloadMuxOut[10] = fifoOut[20][14][w-1];
              unloadMuxOut[11] = fifoOut[21][14][w-1];
              unloadMuxOut[12] = fifoOut[22][14][w-1];
              unloadMuxOut[13] = fifoOut[23][14][w-1];
              unloadMuxOut[14] = fifoOut[24][14][w-1];
              unloadMuxOut[15] = fifoOut[25][14][w-1];
              unloadMuxOut[16] = fifoOut[0][13][w-1];
              unloadMuxOut[17] = fifoOut[1][13][w-1];
              unloadMuxOut[18] = fifoOut[2][13][w-1];
              unloadMuxOut[19] = fifoOut[3][13][w-1];
              unloadMuxOut[20] = fifoOut[4][13][w-1];
              unloadMuxOut[21] = fifoOut[5][13][w-1];
              unloadMuxOut[22] = fifoOut[6][13][w-1];
              unloadMuxOut[23] = fifoOut[7][13][w-1];
              unloadMuxOut[24] = fifoOut[8][13][w-1];
              unloadMuxOut[25] = fifoOut[9][13][w-1];
              unloadMuxOut[26] = fifoOut[10][13][w-1];
              unloadMuxOut[27] = fifoOut[11][13][w-1];
              unloadMuxOut[28] = fifoOut[12][13][w-1];
              unloadMuxOut[29] = fifoOut[13][13][w-1];
              unloadMuxOut[30] = fifoOut[14][13][w-1];
              unloadMuxOut[31] = fifoOut[15][13][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[16][14][w-1];
              unloadMuxOut[1] = fifoOut[17][14][w-1];
              unloadMuxOut[2] = fifoOut[18][14][w-1];
              unloadMuxOut[3] = fifoOut[19][14][w-1];
              unloadMuxOut[4] = fifoOut[20][14][w-1];
              unloadMuxOut[5] = fifoOut[21][14][w-1];
              unloadMuxOut[6] = fifoOut[22][14][w-1];
              unloadMuxOut[7] = fifoOut[23][14][w-1];
              unloadMuxOut[8] = fifoOut[24][14][w-1];
              unloadMuxOut[9] = fifoOut[25][14][w-1];
              unloadMuxOut[10] = fifoOut[0][13][w-1];
              unloadMuxOut[11] = fifoOut[1][13][w-1];
              unloadMuxOut[12] = fifoOut[2][13][w-1];
              unloadMuxOut[13] = fifoOut[3][13][w-1];
              unloadMuxOut[14] = fifoOut[4][13][w-1];
              unloadMuxOut[15] = fifoOut[5][13][w-1];
              unloadMuxOut[16] = fifoOut[6][13][w-1];
              unloadMuxOut[17] = fifoOut[7][13][w-1];
              unloadMuxOut[18] = fifoOut[8][13][w-1];
              unloadMuxOut[19] = fifoOut[9][13][w-1];
              unloadMuxOut[20] = fifoOut[10][13][w-1];
              unloadMuxOut[21] = fifoOut[11][13][w-1];
              unloadMuxOut[22] = fifoOut[12][13][w-1];
              unloadMuxOut[23] = fifoOut[13][13][w-1];
              unloadMuxOut[24] = fifoOut[14][13][w-1];
              unloadMuxOut[25] = fifoOut[15][13][w-1];
              unloadMuxOut[26] = fifoOut[16][13][w-1];
              unloadMuxOut[27] = fifoOut[17][13][w-1];
              unloadMuxOut[28] = fifoOut[18][13][w-1];
              unloadMuxOut[29] = fifoOut[19][13][w-1];
              unloadMuxOut[30] = fifoOut[20][13][w-1];
              unloadMuxOut[31] = fifoOut[21][13][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[22][14][w-1];
              unloadMuxOut[1] = fifoOut[23][14][w-1];
              unloadMuxOut[2] = fifoOut[24][14][w-1];
              unloadMuxOut[3] = fifoOut[25][14][w-1];
              unloadMuxOut[4] = fifoOut[0][13][w-1];
              unloadMuxOut[5] = fifoOut[1][13][w-1];
              unloadMuxOut[6] = fifoOut[2][13][w-1];
              unloadMuxOut[7] = fifoOut[3][13][w-1];
              unloadMuxOut[8] = fifoOut[4][13][w-1];
              unloadMuxOut[9] = fifoOut[5][13][w-1];
              unloadMuxOut[10] = fifoOut[6][13][w-1];
              unloadMuxOut[11] = fifoOut[7][13][w-1];
              unloadMuxOut[12] = fifoOut[8][13][w-1];
              unloadMuxOut[13] = fifoOut[9][13][w-1];
              unloadMuxOut[14] = fifoOut[10][13][w-1];
              unloadMuxOut[15] = fifoOut[11][13][w-1];
              unloadMuxOut[16] = fifoOut[12][13][w-1];
              unloadMuxOut[17] = fifoOut[13][13][w-1];
              unloadMuxOut[18] = fifoOut[14][13][w-1];
              unloadMuxOut[19] = fifoOut[15][13][w-1];
              unloadMuxOut[20] = fifoOut[16][13][w-1];
              unloadMuxOut[21] = fifoOut[17][13][w-1];
              unloadMuxOut[22] = fifoOut[18][13][w-1];
              unloadMuxOut[23] = fifoOut[19][13][w-1];
              unloadMuxOut[24] = fifoOut[20][13][w-1];
              unloadMuxOut[25] = fifoOut[21][13][w-1];
              unloadMuxOut[26] = fifoOut[22][13][w-1];
              unloadMuxOut[27] = fifoOut[23][13][w-1];
              unloadMuxOut[28] = fifoOut[24][13][w-1];
              unloadMuxOut[29] = fifoOut[25][13][w-1];
              unloadMuxOut[30] = fifoOut[0][12][w-1];
              unloadMuxOut[31] = fifoOut[1][12][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[2][13][w-1];
              unloadMuxOut[1] = fifoOut[3][13][w-1];
              unloadMuxOut[2] = fifoOut[4][13][w-1];
              unloadMuxOut[3] = fifoOut[5][13][w-1];
              unloadMuxOut[4] = fifoOut[6][13][w-1];
              unloadMuxOut[5] = fifoOut[7][13][w-1];
              unloadMuxOut[6] = fifoOut[8][13][w-1];
              unloadMuxOut[7] = fifoOut[9][13][w-1];
              unloadMuxOut[8] = fifoOut[10][13][w-1];
              unloadMuxOut[9] = fifoOut[11][13][w-1];
              unloadMuxOut[10] = fifoOut[12][13][w-1];
              unloadMuxOut[11] = fifoOut[13][13][w-1];
              unloadMuxOut[12] = fifoOut[14][13][w-1];
              unloadMuxOut[13] = fifoOut[15][13][w-1];
              unloadMuxOut[14] = fifoOut[16][13][w-1];
              unloadMuxOut[15] = fifoOut[17][13][w-1];
              unloadMuxOut[16] = fifoOut[18][13][w-1];
              unloadMuxOut[17] = fifoOut[19][13][w-1];
              unloadMuxOut[18] = fifoOut[20][13][w-1];
              unloadMuxOut[19] = fifoOut[21][13][w-1];
              unloadMuxOut[20] = fifoOut[22][13][w-1];
              unloadMuxOut[21] = fifoOut[23][13][w-1];
              unloadMuxOut[22] = fifoOut[24][13][w-1];
              unloadMuxOut[23] = fifoOut[25][13][w-1];
              unloadMuxOut[24] = fifoOut[0][12][w-1];
              unloadMuxOut[25] = fifoOut[1][12][w-1];
              unloadMuxOut[26] = fifoOut[26][16][w-1];
              unloadMuxOut[27] = fifoOut[27][16][w-1];
              unloadMuxOut[28] = fifoOut[28][16][w-1];
              unloadMuxOut[29] = fifoOut[29][16][w-1];
              unloadMuxOut[30] = fifoOut[30][16][w-1];
              unloadMuxOut[31] = fifoOut[31][16][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[8][13][w-1];
              unloadMuxOut[1] = fifoOut[9][13][w-1];
              unloadMuxOut[2] = fifoOut[10][13][w-1];
              unloadMuxOut[3] = fifoOut[11][13][w-1];
              unloadMuxOut[4] = fifoOut[12][13][w-1];
              unloadMuxOut[5] = fifoOut[13][13][w-1];
              unloadMuxOut[6] = fifoOut[14][13][w-1];
              unloadMuxOut[7] = fifoOut[15][13][w-1];
              unloadMuxOut[8] = fifoOut[16][13][w-1];
              unloadMuxOut[9] = fifoOut[17][13][w-1];
              unloadMuxOut[10] = fifoOut[18][13][w-1];
              unloadMuxOut[11] = fifoOut[19][13][w-1];
              unloadMuxOut[12] = fifoOut[20][13][w-1];
              unloadMuxOut[13] = fifoOut[21][13][w-1];
              unloadMuxOut[14] = fifoOut[22][13][w-1];
              unloadMuxOut[15] = fifoOut[23][13][w-1];
              unloadMuxOut[16] = fifoOut[24][13][w-1];
              unloadMuxOut[17] = fifoOut[25][13][w-1];
              unloadMuxOut[18] = fifoOut[0][12][w-1];
              unloadMuxOut[19] = fifoOut[1][12][w-1];
              unloadMuxOut[20] = fifoOut[26][16][w-1];
              unloadMuxOut[21] = fifoOut[27][16][w-1];
              unloadMuxOut[22] = fifoOut[28][16][w-1];
              unloadMuxOut[23] = fifoOut[29][16][w-1];
              unloadMuxOut[24] = fifoOut[30][16][w-1];
              unloadMuxOut[25] = fifoOut[31][16][w-1];
              unloadMuxOut[26] = fifoOut[32][16][w-1];
              unloadMuxOut[27] = fifoOut[33][16][w-1];
              unloadMuxOut[28] = fifoOut[34][16][w-1];
              unloadMuxOut[29] = fifoOut[35][16][w-1];
              unloadMuxOut[30] = fifoOut[36][16][w-1];
              unloadMuxOut[31] = fifoOut[37][16][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[14][13][w-1];
              unloadMuxOut[1] = fifoOut[15][13][w-1];
              unloadMuxOut[2] = fifoOut[16][13][w-1];
              unloadMuxOut[3] = fifoOut[17][13][w-1];
              unloadMuxOut[4] = fifoOut[18][13][w-1];
              unloadMuxOut[5] = fifoOut[19][13][w-1];
              unloadMuxOut[6] = fifoOut[20][13][w-1];
              unloadMuxOut[7] = fifoOut[21][13][w-1];
              unloadMuxOut[8] = fifoOut[22][13][w-1];
              unloadMuxOut[9] = fifoOut[23][13][w-1];
              unloadMuxOut[10] = fifoOut[24][13][w-1];
              unloadMuxOut[11] = fifoOut[25][13][w-1];
              unloadMuxOut[12] = fifoOut[0][12][w-1];
              unloadMuxOut[13] = fifoOut[1][12][w-1];
              unloadMuxOut[14] = fifoOut[26][16][w-1];
              unloadMuxOut[15] = fifoOut[27][16][w-1];
              unloadMuxOut[16] = fifoOut[28][16][w-1];
              unloadMuxOut[17] = fifoOut[29][16][w-1];
              unloadMuxOut[18] = fifoOut[30][16][w-1];
              unloadMuxOut[19] = fifoOut[31][16][w-1];
              unloadMuxOut[20] = fifoOut[32][16][w-1];
              unloadMuxOut[21] = fifoOut[33][16][w-1];
              unloadMuxOut[22] = fifoOut[34][16][w-1];
              unloadMuxOut[23] = fifoOut[35][16][w-1];
              unloadMuxOut[24] = fifoOut[36][16][w-1];
              unloadMuxOut[25] = fifoOut[37][16][w-1];
              unloadMuxOut[26] = fifoOut[38][16][w-1];
              unloadMuxOut[27] = fifoOut[39][16][w-1];
              unloadMuxOut[28] = fifoOut[40][16][w-1];
              unloadMuxOut[29] = fifoOut[41][16][w-1];
              unloadMuxOut[30] = fifoOut[42][16][w-1];
              unloadMuxOut[31] = fifoOut[43][16][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[20][13][w-1];
              unloadMuxOut[1] = fifoOut[21][13][w-1];
              unloadMuxOut[2] = fifoOut[22][13][w-1];
              unloadMuxOut[3] = fifoOut[23][13][w-1];
              unloadMuxOut[4] = fifoOut[24][13][w-1];
              unloadMuxOut[5] = fifoOut[25][13][w-1];
              unloadMuxOut[6] = fifoOut[0][12][w-1];
              unloadMuxOut[7] = fifoOut[1][12][w-1];
              unloadMuxOut[8] = fifoOut[26][16][w-1];
              unloadMuxOut[9] = fifoOut[27][16][w-1];
              unloadMuxOut[10] = fifoOut[28][16][w-1];
              unloadMuxOut[11] = fifoOut[29][16][w-1];
              unloadMuxOut[12] = fifoOut[30][16][w-1];
              unloadMuxOut[13] = fifoOut[31][16][w-1];
              unloadMuxOut[14] = fifoOut[32][16][w-1];
              unloadMuxOut[15] = fifoOut[33][16][w-1];
              unloadMuxOut[16] = fifoOut[34][16][w-1];
              unloadMuxOut[17] = fifoOut[35][16][w-1];
              unloadMuxOut[18] = fifoOut[36][16][w-1];
              unloadMuxOut[19] = fifoOut[37][16][w-1];
              unloadMuxOut[20] = fifoOut[38][16][w-1];
              unloadMuxOut[21] = fifoOut[39][16][w-1];
              unloadMuxOut[22] = fifoOut[40][16][w-1];
              unloadMuxOut[23] = fifoOut[41][16][w-1];
              unloadMuxOut[24] = fifoOut[42][16][w-1];
              unloadMuxOut[25] = fifoOut[43][16][w-1];
              unloadMuxOut[26] = fifoOut[44][16][w-1];
              unloadMuxOut[27] = fifoOut[45][16][w-1];
              unloadMuxOut[28] = fifoOut[46][16][w-1];
              unloadMuxOut[29] = fifoOut[47][16][w-1];
              unloadMuxOut[30] = fifoOut[48][16][w-1];
              unloadMuxOut[31] = fifoOut[49][16][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[0][12][w-1];
              unloadMuxOut[1] = fifoOut[1][12][w-1];
              unloadMuxOut[2] = fifoOut[26][16][w-1];
              unloadMuxOut[3] = fifoOut[27][16][w-1];
              unloadMuxOut[4] = fifoOut[28][16][w-1];
              unloadMuxOut[5] = fifoOut[29][16][w-1];
              unloadMuxOut[6] = fifoOut[30][16][w-1];
              unloadMuxOut[7] = fifoOut[31][16][w-1];
              unloadMuxOut[8] = fifoOut[32][16][w-1];
              unloadMuxOut[9] = fifoOut[33][16][w-1];
              unloadMuxOut[10] = fifoOut[34][16][w-1];
              unloadMuxOut[11] = fifoOut[35][16][w-1];
              unloadMuxOut[12] = fifoOut[36][16][w-1];
              unloadMuxOut[13] = fifoOut[37][16][w-1];
              unloadMuxOut[14] = fifoOut[38][16][w-1];
              unloadMuxOut[15] = fifoOut[39][16][w-1];
              unloadMuxOut[16] = fifoOut[40][16][w-1];
              unloadMuxOut[17] = fifoOut[41][16][w-1];
              unloadMuxOut[18] = fifoOut[42][16][w-1];
              unloadMuxOut[19] = fifoOut[43][16][w-1];
              unloadMuxOut[20] = fifoOut[44][16][w-1];
              unloadMuxOut[21] = fifoOut[45][16][w-1];
              unloadMuxOut[22] = fifoOut[46][16][w-1];
              unloadMuxOut[23] = fifoOut[47][16][w-1];
              unloadMuxOut[24] = fifoOut[48][16][w-1];
              unloadMuxOut[25] = fifoOut[49][16][w-1];
              unloadMuxOut[26] = fifoOut[50][16][w-1];
              unloadMuxOut[27] = fifoOut[51][16][w-1];
              unloadMuxOut[28] = fifoOut[26][15][w-1];
              unloadMuxOut[29] = fifoOut[27][15][w-1];
              unloadMuxOut[30] = fifoOut[28][15][w-1];
              unloadMuxOut[31] = fifoOut[29][15][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[30][16][w-1];
              unloadMuxOut[1] = fifoOut[31][16][w-1];
              unloadMuxOut[2] = fifoOut[32][16][w-1];
              unloadMuxOut[3] = fifoOut[33][16][w-1];
              unloadMuxOut[4] = fifoOut[34][16][w-1];
              unloadMuxOut[5] = fifoOut[35][16][w-1];
              unloadMuxOut[6] = fifoOut[36][16][w-1];
              unloadMuxOut[7] = fifoOut[37][16][w-1];
              unloadMuxOut[8] = fifoOut[38][16][w-1];
              unloadMuxOut[9] = fifoOut[39][16][w-1];
              unloadMuxOut[10] = fifoOut[40][16][w-1];
              unloadMuxOut[11] = fifoOut[41][16][w-1];
              unloadMuxOut[12] = fifoOut[42][16][w-1];
              unloadMuxOut[13] = fifoOut[43][16][w-1];
              unloadMuxOut[14] = fifoOut[44][16][w-1];
              unloadMuxOut[15] = fifoOut[45][16][w-1];
              unloadMuxOut[16] = fifoOut[46][16][w-1];
              unloadMuxOut[17] = fifoOut[47][16][w-1];
              unloadMuxOut[18] = fifoOut[48][16][w-1];
              unloadMuxOut[19] = fifoOut[49][16][w-1];
              unloadMuxOut[20] = fifoOut[50][16][w-1];
              unloadMuxOut[21] = fifoOut[51][16][w-1];
              unloadMuxOut[22] = fifoOut[26][15][w-1];
              unloadMuxOut[23] = fifoOut[27][15][w-1];
              unloadMuxOut[24] = fifoOut[28][15][w-1];
              unloadMuxOut[25] = fifoOut[29][15][w-1];
              unloadMuxOut[26] = fifoOut[30][15][w-1];
              unloadMuxOut[27] = fifoOut[31][15][w-1];
              unloadMuxOut[28] = fifoOut[32][15][w-1];
              unloadMuxOut[29] = fifoOut[33][15][w-1];
              unloadMuxOut[30] = fifoOut[34][15][w-1];
              unloadMuxOut[31] = fifoOut[35][15][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[36][16][w-1];
              unloadMuxOut[1] = fifoOut[37][16][w-1];
              unloadMuxOut[2] = fifoOut[38][16][w-1];
              unloadMuxOut[3] = fifoOut[39][16][w-1];
              unloadMuxOut[4] = fifoOut[40][16][w-1];
              unloadMuxOut[5] = fifoOut[41][16][w-1];
              unloadMuxOut[6] = fifoOut[42][16][w-1];
              unloadMuxOut[7] = fifoOut[43][16][w-1];
              unloadMuxOut[8] = fifoOut[44][16][w-1];
              unloadMuxOut[9] = fifoOut[45][16][w-1];
              unloadMuxOut[10] = fifoOut[46][16][w-1];
              unloadMuxOut[11] = fifoOut[47][16][w-1];
              unloadMuxOut[12] = fifoOut[48][16][w-1];
              unloadMuxOut[13] = fifoOut[49][16][w-1];
              unloadMuxOut[14] = fifoOut[50][16][w-1];
              unloadMuxOut[15] = fifoOut[51][16][w-1];
              unloadMuxOut[16] = fifoOut[26][15][w-1];
              unloadMuxOut[17] = fifoOut[27][15][w-1];
              unloadMuxOut[18] = fifoOut[28][15][w-1];
              unloadMuxOut[19] = fifoOut[29][15][w-1];
              unloadMuxOut[20] = fifoOut[30][15][w-1];
              unloadMuxOut[21] = fifoOut[31][15][w-1];
              unloadMuxOut[22] = fifoOut[32][15][w-1];
              unloadMuxOut[23] = fifoOut[33][15][w-1];
              unloadMuxOut[24] = fifoOut[34][15][w-1];
              unloadMuxOut[25] = fifoOut[35][15][w-1];
              unloadMuxOut[26] = fifoOut[36][15][w-1];
              unloadMuxOut[27] = fifoOut[37][15][w-1];
              unloadMuxOut[28] = fifoOut[38][15][w-1];
              unloadMuxOut[29] = fifoOut[39][15][w-1];
              unloadMuxOut[30] = fifoOut[40][15][w-1];
              unloadMuxOut[31] = fifoOut[41][15][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[42][16][w-1];
              unloadMuxOut[1] = fifoOut[43][16][w-1];
              unloadMuxOut[2] = fifoOut[44][16][w-1];
              unloadMuxOut[3] = fifoOut[45][16][w-1];
              unloadMuxOut[4] = fifoOut[46][16][w-1];
              unloadMuxOut[5] = fifoOut[47][16][w-1];
              unloadMuxOut[6] = fifoOut[48][16][w-1];
              unloadMuxOut[7] = fifoOut[49][16][w-1];
              unloadMuxOut[8] = fifoOut[50][16][w-1];
              unloadMuxOut[9] = fifoOut[51][16][w-1];
              unloadMuxOut[10] = fifoOut[26][15][w-1];
              unloadMuxOut[11] = fifoOut[27][15][w-1];
              unloadMuxOut[12] = fifoOut[28][15][w-1];
              unloadMuxOut[13] = fifoOut[29][15][w-1];
              unloadMuxOut[14] = fifoOut[30][15][w-1];
              unloadMuxOut[15] = fifoOut[31][15][w-1];
              unloadMuxOut[16] = fifoOut[32][15][w-1];
              unloadMuxOut[17] = fifoOut[33][15][w-1];
              unloadMuxOut[18] = fifoOut[34][15][w-1];
              unloadMuxOut[19] = fifoOut[35][15][w-1];
              unloadMuxOut[20] = fifoOut[36][15][w-1];
              unloadMuxOut[21] = fifoOut[37][15][w-1];
              unloadMuxOut[22] = fifoOut[38][15][w-1];
              unloadMuxOut[23] = fifoOut[39][15][w-1];
              unloadMuxOut[24] = fifoOut[40][15][w-1];
              unloadMuxOut[25] = fifoOut[41][15][w-1];
              unloadMuxOut[26] = fifoOut[42][15][w-1];
              unloadMuxOut[27] = fifoOut[43][15][w-1];
              unloadMuxOut[28] = fifoOut[44][15][w-1];
              unloadMuxOut[29] = fifoOut[45][15][w-1];
              unloadMuxOut[30] = fifoOut[46][15][w-1];
              unloadMuxOut[31] = fifoOut[47][15][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[48][16][w-1];
              unloadMuxOut[1] = fifoOut[49][16][w-1];
              unloadMuxOut[2] = fifoOut[50][16][w-1];
              unloadMuxOut[3] = fifoOut[51][16][w-1];
              unloadMuxOut[4] = fifoOut[26][15][w-1];
              unloadMuxOut[5] = fifoOut[27][15][w-1];
              unloadMuxOut[6] = fifoOut[28][15][w-1];
              unloadMuxOut[7] = fifoOut[29][15][w-1];
              unloadMuxOut[8] = fifoOut[30][15][w-1];
              unloadMuxOut[9] = fifoOut[31][15][w-1];
              unloadMuxOut[10] = fifoOut[32][15][w-1];
              unloadMuxOut[11] = fifoOut[33][15][w-1];
              unloadMuxOut[12] = fifoOut[34][15][w-1];
              unloadMuxOut[13] = fifoOut[35][15][w-1];
              unloadMuxOut[14] = fifoOut[36][15][w-1];
              unloadMuxOut[15] = fifoOut[37][15][w-1];
              unloadMuxOut[16] = fifoOut[38][15][w-1];
              unloadMuxOut[17] = fifoOut[39][15][w-1];
              unloadMuxOut[18] = fifoOut[40][15][w-1];
              unloadMuxOut[19] = fifoOut[41][15][w-1];
              unloadMuxOut[20] = fifoOut[42][15][w-1];
              unloadMuxOut[21] = fifoOut[43][15][w-1];
              unloadMuxOut[22] = fifoOut[44][15][w-1];
              unloadMuxOut[23] = fifoOut[45][15][w-1];
              unloadMuxOut[24] = fifoOut[46][15][w-1];
              unloadMuxOut[25] = fifoOut[47][15][w-1];
              unloadMuxOut[26] = fifoOut[48][15][w-1];
              unloadMuxOut[27] = fifoOut[49][15][w-1];
              unloadMuxOut[28] = fifoOut[50][15][w-1];
              unloadMuxOut[29] = fifoOut[51][15][w-1];
              unloadMuxOut[30] = fifoOut[26][14][w-1];
              unloadMuxOut[31] = fifoOut[27][14][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[28][15][w-1];
              unloadMuxOut[1] = fifoOut[29][15][w-1];
              unloadMuxOut[2] = fifoOut[30][15][w-1];
              unloadMuxOut[3] = fifoOut[31][15][w-1];
              unloadMuxOut[4] = fifoOut[32][15][w-1];
              unloadMuxOut[5] = fifoOut[33][15][w-1];
              unloadMuxOut[6] = fifoOut[34][15][w-1];
              unloadMuxOut[7] = fifoOut[35][15][w-1];
              unloadMuxOut[8] = fifoOut[36][15][w-1];
              unloadMuxOut[9] = fifoOut[37][15][w-1];
              unloadMuxOut[10] = fifoOut[38][15][w-1];
              unloadMuxOut[11] = fifoOut[39][15][w-1];
              unloadMuxOut[12] = fifoOut[40][15][w-1];
              unloadMuxOut[13] = fifoOut[41][15][w-1];
              unloadMuxOut[14] = fifoOut[42][15][w-1];
              unloadMuxOut[15] = fifoOut[43][15][w-1];
              unloadMuxOut[16] = fifoOut[44][15][w-1];
              unloadMuxOut[17] = fifoOut[45][15][w-1];
              unloadMuxOut[18] = fifoOut[46][15][w-1];
              unloadMuxOut[19] = fifoOut[47][15][w-1];
              unloadMuxOut[20] = fifoOut[48][15][w-1];
              unloadMuxOut[21] = fifoOut[49][15][w-1];
              unloadMuxOut[22] = fifoOut[50][15][w-1];
              unloadMuxOut[23] = fifoOut[51][15][w-1];
              unloadMuxOut[24] = fifoOut[26][14][w-1];
              unloadMuxOut[25] = fifoOut[27][14][w-1];
              unloadMuxOut[26] = fifoOut[28][14][w-1];
              unloadMuxOut[27] = fifoOut[29][14][w-1];
              unloadMuxOut[28] = fifoOut[30][14][w-1];
              unloadMuxOut[29] = fifoOut[31][14][w-1];
              unloadMuxOut[30] = fifoOut[32][14][w-1];
              unloadMuxOut[31] = fifoOut[33][14][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[34][15][w-1];
              unloadMuxOut[1] = fifoOut[35][15][w-1];
              unloadMuxOut[2] = fifoOut[36][15][w-1];
              unloadMuxOut[3] = fifoOut[37][15][w-1];
              unloadMuxOut[4] = fifoOut[38][15][w-1];
              unloadMuxOut[5] = fifoOut[39][15][w-1];
              unloadMuxOut[6] = fifoOut[40][15][w-1];
              unloadMuxOut[7] = fifoOut[41][15][w-1];
              unloadMuxOut[8] = fifoOut[42][15][w-1];
              unloadMuxOut[9] = fifoOut[2][13][w-1];
              unloadMuxOut[10] = fifoOut[3][13][w-1];
              unloadMuxOut[11] = fifoOut[4][13][w-1];
              unloadMuxOut[12] = fifoOut[5][13][w-1];
              unloadMuxOut[13] = fifoOut[6][13][w-1];
              unloadMuxOut[14] = fifoOut[7][13][w-1];
              unloadMuxOut[15] = fifoOut[8][13][w-1];
              unloadMuxOut[16] = fifoOut[9][13][w-1];
              unloadMuxOut[17] = fifoOut[10][13][w-1];
              unloadMuxOut[18] = fifoOut[11][13][w-1];
              unloadMuxOut[19] = fifoOut[12][13][w-1];
              unloadMuxOut[20] = fifoOut[13][13][w-1];
              unloadMuxOut[21] = fifoOut[14][13][w-1];
              unloadMuxOut[22] = fifoOut[15][13][w-1];
              unloadMuxOut[23] = fifoOut[16][13][w-1];
              unloadMuxOut[24] = fifoOut[17][13][w-1];
              unloadMuxOut[25] = fifoOut[18][13][w-1];
              unloadMuxOut[26] = fifoOut[19][13][w-1];
              unloadMuxOut[27] = fifoOut[20][13][w-1];
              unloadMuxOut[28] = fifoOut[21][13][w-1];
              unloadMuxOut[29] = fifoOut[22][13][w-1];
              unloadMuxOut[30] = fifoOut[23][13][w-1];
              unloadMuxOut[31] = fifoOut[24][13][w-1];
       end
       16: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0; 
             end
       end
    endcase //unload case end
    case(iteration_0_indicator)
       0: begin
         case(rd_address_case)
         0: begin
              muxOutConnector[0] = fifoOut[35][10];
              muxOutConnector[1] = fifoOut[36][10];
              muxOutConnector[2] = fifoOut[37][10];
              muxOutConnector[3] = fifoOut[38][10];
              muxOutConnector[4] = fifoOut[39][10];
              muxOutConnector[5] = fifoOut[40][10];
              muxOutConnector[6] = fifoOut[41][10];
              muxOutConnector[7] = fifoOut[42][10];
              muxOutConnector[8] = fifoOut[43][10];
              muxOutConnector[9] = fifoOut[44][10];
              muxOutConnector[10] = fifoOut[45][10];
              muxOutConnector[11] = fifoOut[46][10];
              muxOutConnector[12] = fifoOut[47][10];
              muxOutConnector[13] = fifoOut[48][10];
              muxOutConnector[14] = fifoOut[49][10];
              muxOutConnector[15] = fifoOut[50][10];
              muxOutConnector[16] = fifoOut[51][10];
              muxOutConnector[17] = fifoOut[26][9];
              muxOutConnector[18] = fifoOut[27][9];
              muxOutConnector[19] = fifoOut[28][9];
              muxOutConnector[20] = fifoOut[29][9];
              muxOutConnector[21] = fifoOut[30][9];
              muxOutConnector[22] = fifoOut[31][9];
              muxOutConnector[23] = fifoOut[32][9];
              muxOutConnector[24] = fifoOut[33][9];
              muxOutConnector[25] = fifoOut[34][9];
              muxOutConnector[26] = fifoOut[30][0];
              muxOutConnector[27] = fifoOut[31][0];
              muxOutConnector[28] = fifoOut[32][0];
              muxOutConnector[29] = fifoOut[33][0];
              muxOutConnector[30] = fifoOut[34][0];
              muxOutConnector[31] = fifoOut[35][0];
              muxOutConnector[32] = fifoOut[36][0];
              muxOutConnector[33] = fifoOut[37][0];
              muxOutConnector[34] = fifoOut[38][0];
              muxOutConnector[35] = fifoOut[39][0];
              muxOutConnector[36] = fifoOut[40][0];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         1: begin
              muxOutConnector[0] = fifoOut[35][10];
              muxOutConnector[1] = fifoOut[36][10];
              muxOutConnector[2] = fifoOut[37][10];
              muxOutConnector[3] = fifoOut[38][10];
              muxOutConnector[4] = fifoOut[39][10];
              muxOutConnector[5] = fifoOut[40][10];
              muxOutConnector[6] = fifoOut[41][10];
              muxOutConnector[7] = fifoOut[42][10];
              muxOutConnector[8] = fifoOut[43][10];
              muxOutConnector[9] = fifoOut[44][10];
              muxOutConnector[10] = fifoOut[45][10];
              muxOutConnector[11] = fifoOut[46][10];
              muxOutConnector[12] = fifoOut[47][10];
              muxOutConnector[13] = fifoOut[48][10];
              muxOutConnector[14] = fifoOut[49][10];
              muxOutConnector[15] = fifoOut[50][10];
              muxOutConnector[16] = fifoOut[51][10];
              muxOutConnector[17] = fifoOut[26][9];
              muxOutConnector[18] = fifoOut[27][9];
              muxOutConnector[19] = fifoOut[28][9];
              muxOutConnector[20] = fifoOut[29][9];
              muxOutConnector[21] = fifoOut[30][9];
              muxOutConnector[22] = fifoOut[31][9];
              muxOutConnector[23] = fifoOut[32][9];
              muxOutConnector[24] = fifoOut[33][9];
              muxOutConnector[25] = fifoOut[34][9];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         2: begin
              muxOutConnector[0] = fifoOut[35][10];
              muxOutConnector[1] = fifoOut[36][10];
              muxOutConnector[2] = fifoOut[37][10];
              muxOutConnector[3] = fifoOut[38][10];
              muxOutConnector[4] = fifoOut[39][10];
              muxOutConnector[5] = fifoOut[40][10];
              muxOutConnector[6] = fifoOut[41][10];
              muxOutConnector[7] = fifoOut[42][10];
              muxOutConnector[8] = fifoOut[43][10];
              muxOutConnector[9] = fifoOut[44][10];
              muxOutConnector[10] = fifoOut[45][10];
              muxOutConnector[11] = fifoOut[46][10];
              muxOutConnector[12] = fifoOut[47][10];
              muxOutConnector[13] = fifoOut[48][10];
              muxOutConnector[14] = fifoOut[49][10];
              muxOutConnector[15] = fifoOut[50][10];
              muxOutConnector[16] = fifoOut[51][10];
              muxOutConnector[17] = fifoOut[26][9];
              muxOutConnector[18] = fifoOut[27][9];
              muxOutConnector[19] = fifoOut[28][9];
              muxOutConnector[20] = fifoOut[29][9];
              muxOutConnector[21] = fifoOut[30][9];
              muxOutConnector[22] = fifoOut[31][9];
              muxOutConnector[23] = fifoOut[32][9];
              muxOutConnector[24] = fifoOut[33][9];
              muxOutConnector[25] = fifoOut[34][9];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         3: begin
              muxOutConnector[0] = fifoOut[35][10];
              muxOutConnector[1] = fifoOut[36][10];
              muxOutConnector[2] = fifoOut[37][10];
              muxOutConnector[3] = fifoOut[38][10];
              muxOutConnector[4] = fifoOut[39][10];
              muxOutConnector[5] = fifoOut[40][10];
              muxOutConnector[6] = fifoOut[41][10];
              muxOutConnector[7] = fifoOut[42][10];
              muxOutConnector[8] = fifoOut[43][10];
              muxOutConnector[9] = fifoOut[44][10];
              muxOutConnector[10] = fifoOut[45][10];
              muxOutConnector[11] = fifoOut[46][10];
              muxOutConnector[12] = fifoOut[47][10];
              muxOutConnector[13] = fifoOut[48][10];
              muxOutConnector[14] = fifoOut[49][10];
              muxOutConnector[15] = fifoOut[50][10];
              muxOutConnector[16] = fifoOut[51][10];
              muxOutConnector[17] = fifoOut[26][9];
              muxOutConnector[18] = fifoOut[27][9];
              muxOutConnector[19] = fifoOut[28][9];
              muxOutConnector[20] = fifoOut[29][9];
              muxOutConnector[21] = fifoOut[30][9];
              muxOutConnector[22] = fifoOut[31][9];
              muxOutConnector[23] = fifoOut[32][9];
              muxOutConnector[24] = fifoOut[33][9];
              muxOutConnector[25] = fifoOut[34][9];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         4: begin
              muxOutConnector[0] = fifoOut[35][10];
              muxOutConnector[1] = fifoOut[36][10];
              muxOutConnector[2] = fifoOut[37][10];
              muxOutConnector[3] = fifoOut[38][10];
              muxOutConnector[4] = fifoOut[39][10];
              muxOutConnector[5] = fifoOut[40][10];
              muxOutConnector[6] = fifoOut[41][10];
              muxOutConnector[7] = fifoOut[42][10];
              muxOutConnector[8] = fifoOut[43][10];
              muxOutConnector[9] = fifoOut[44][10];
              muxOutConnector[10] = fifoOut[45][10];
              muxOutConnector[11] = fifoOut[46][10];
              muxOutConnector[12] = fifoOut[47][10];
              muxOutConnector[13] = fifoOut[48][10];
              muxOutConnector[14] = fifoOut[49][10];
              muxOutConnector[15] = fifoOut[50][10];
              muxOutConnector[16] = fifoOut[51][10];
              muxOutConnector[17] = fifoOut[26][9];
              muxOutConnector[18] = fifoOut[27][9];
              muxOutConnector[19] = fifoOut[28][9];
              muxOutConnector[20] = fifoOut[29][9];
              muxOutConnector[21] = fifoOut[30][9];
              muxOutConnector[22] = fifoOut[31][9];
              muxOutConnector[23] = fifoOut[32][9];
              muxOutConnector[24] = fifoOut[33][9];
              muxOutConnector[25] = fifoOut[34][9];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         5: begin
              muxOutConnector[0] = fifoOut[35][10];
              muxOutConnector[1] = fifoOut[36][10];
              muxOutConnector[2] = fifoOut[37][10];
              muxOutConnector[3] = fifoOut[38][10];
              muxOutConnector[4] = fifoOut[39][10];
              muxOutConnector[5] = fifoOut[40][10];
              muxOutConnector[6] = fifoOut[41][10];
              muxOutConnector[7] = fifoOut[42][10];
              muxOutConnector[8] = fifoOut[43][10];
              muxOutConnector[9] = fifoOut[44][10];
              muxOutConnector[10] = fifoOut[45][10];
              muxOutConnector[11] = fifoOut[46][10];
              muxOutConnector[12] = fifoOut[47][10];
              muxOutConnector[13] = fifoOut[48][10];
              muxOutConnector[14] = fifoOut[49][10];
              muxOutConnector[15] = fifoOut[50][10];
              muxOutConnector[16] = fifoOut[51][10];
              muxOutConnector[17] = fifoOut[26][9];
              muxOutConnector[18] = fifoOut[27][9];
              muxOutConnector[19] = fifoOut[28][9];
              muxOutConnector[20] = fifoOut[29][9];
              muxOutConnector[21] = fifoOut[30][9];
              muxOutConnector[22] = fifoOut[31][9];
              muxOutConnector[23] = fifoOut[32][9];
              muxOutConnector[24] = fifoOut[33][9];
              muxOutConnector[25] = fifoOut[34][9];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         6: begin
              muxOutConnector[0] = fifoOut[35][10];
              muxOutConnector[1] = fifoOut[36][10];
              muxOutConnector[2] = fifoOut[37][10];
              muxOutConnector[3] = fifoOut[38][10];
              muxOutConnector[4] = fifoOut[39][10];
              muxOutConnector[5] = fifoOut[40][10];
              muxOutConnector[6] = fifoOut[41][10];
              muxOutConnector[7] = fifoOut[42][10];
              muxOutConnector[8] = fifoOut[43][10];
              muxOutConnector[9] = fifoOut[44][10];
              muxOutConnector[10] = fifoOut[45][10];
              muxOutConnector[11] = fifoOut[46][10];
              muxOutConnector[12] = fifoOut[47][10];
              muxOutConnector[13] = fifoOut[48][10];
              muxOutConnector[14] = fifoOut[49][10];
              muxOutConnector[15] = fifoOut[50][10];
              muxOutConnector[16] = fifoOut[51][10];
              muxOutConnector[17] = fifoOut[26][9];
              muxOutConnector[18] = fifoOut[27][9];
              muxOutConnector[19] = fifoOut[28][9];
              muxOutConnector[20] = fifoOut[29][9];
              muxOutConnector[21] = fifoOut[30][9];
              muxOutConnector[22] = fifoOut[31][9];
              muxOutConnector[23] = fifoOut[32][9];
              muxOutConnector[24] = fifoOut[33][9];
              muxOutConnector[25] = fifoOut[34][9];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         7: begin
              muxOutConnector[0] = fifoOut[35][10];
              muxOutConnector[1] = fifoOut[36][10];
              muxOutConnector[2] = fifoOut[37][10];
              muxOutConnector[3] = fifoOut[38][10];
              muxOutConnector[4] = fifoOut[39][10];
              muxOutConnector[5] = fifoOut[40][10];
              muxOutConnector[6] = fifoOut[41][10];
              muxOutConnector[7] = fifoOut[42][10];
              muxOutConnector[8] = fifoOut[43][10];
              muxOutConnector[9] = fifoOut[44][10];
              muxOutConnector[10] = fifoOut[45][10];
              muxOutConnector[11] = fifoOut[46][10];
              muxOutConnector[12] = fifoOut[47][10];
              muxOutConnector[13] = fifoOut[48][10];
              muxOutConnector[14] = fifoOut[49][10];
              muxOutConnector[15] = fifoOut[50][10];
              muxOutConnector[16] = fifoOut[51][10];
              muxOutConnector[17] = fifoOut[26][9];
              muxOutConnector[18] = fifoOut[27][9];
              muxOutConnector[19] = fifoOut[28][9];
              muxOutConnector[20] = fifoOut[29][9];
              muxOutConnector[21] = fifoOut[30][9];
              muxOutConnector[22] = fifoOut[31][9];
              muxOutConnector[23] = fifoOut[32][9];
              muxOutConnector[24] = fifoOut[33][9];
              muxOutConnector[25] = fifoOut[34][9];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         8: begin
              muxOutConnector[0] = fifoOut[35][10];
              muxOutConnector[1] = fifoOut[36][10];
              muxOutConnector[2] = fifoOut[37][10];
              muxOutConnector[3] = fifoOut[38][10];
              muxOutConnector[4] = fifoOut[39][10];
              muxOutConnector[5] = fifoOut[40][10];
              muxOutConnector[6] = fifoOut[41][10];
              muxOutConnector[7] = fifoOut[42][10];
              muxOutConnector[8] = fifoOut[43][10];
              muxOutConnector[9] = fifoOut[44][10];
              muxOutConnector[10] = fifoOut[45][10];
              muxOutConnector[11] = fifoOut[46][10];
              muxOutConnector[12] = fifoOut[47][10];
              muxOutConnector[13] = fifoOut[48][10];
              muxOutConnector[14] = fifoOut[49][10];
              muxOutConnector[15] = fifoOut[50][10];
              muxOutConnector[16] = fifoOut[51][10];
              muxOutConnector[17] = fifoOut[26][9];
              muxOutConnector[18] = fifoOut[27][9];
              muxOutConnector[19] = fifoOut[28][9];
              muxOutConnector[20] = fifoOut[29][9];
              muxOutConnector[21] = fifoOut[30][9];
              muxOutConnector[22] = fifoOut[31][9];
              muxOutConnector[23] = fifoOut[32][9];
              muxOutConnector[24] = fifoOut[33][9];
              muxOutConnector[25] = fifoOut[34][9];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         9: begin
              muxOutConnector[0] = fifoOut[35][10];
              muxOutConnector[1] = fifoOut[36][10];
              muxOutConnector[2] = fifoOut[37][10];
              muxOutConnector[3] = fifoOut[38][10];
              muxOutConnector[4] = fifoOut[39][10];
              muxOutConnector[5] = fifoOut[40][10];
              muxOutConnector[6] = fifoOut[41][10];
              muxOutConnector[7] = fifoOut[42][10];
              muxOutConnector[8] = fifoOut[43][10];
              muxOutConnector[9] = fifoOut[44][10];
              muxOutConnector[10] = fifoOut[45][10];
              muxOutConnector[11] = fifoOut[46][10];
              muxOutConnector[12] = fifoOut[47][10];
              muxOutConnector[13] = fifoOut[48][10];
              muxOutConnector[14] = fifoOut[49][10];
              muxOutConnector[15] = fifoOut[50][10];
              muxOutConnector[16] = fifoOut[51][10];
              muxOutConnector[17] = fifoOut[26][9];
              muxOutConnector[18] = fifoOut[27][9];
              muxOutConnector[19] = fifoOut[28][9];
              muxOutConnector[20] = fifoOut[29][9];
              muxOutConnector[21] = fifoOut[30][9];
              muxOutConnector[22] = fifoOut[31][9];
              muxOutConnector[23] = fifoOut[32][9];
              muxOutConnector[24] = fifoOut[33][9];
              muxOutConnector[25] = fifoOut[34][9];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         10: begin
              muxOutConnector[0] = fifoOut[35][10];
              muxOutConnector[1] = fifoOut[36][10];
              muxOutConnector[2] = fifoOut[37][10];
              muxOutConnector[3] = fifoOut[38][10];
              muxOutConnector[4] = fifoOut[39][10];
              muxOutConnector[5] = fifoOut[40][10];
              muxOutConnector[6] = fifoOut[41][10];
              muxOutConnector[7] = fifoOut[42][10];
              muxOutConnector[8] = fifoOut[2][8];
              muxOutConnector[9] = fifoOut[3][8];
              muxOutConnector[10] = fifoOut[4][8];
              muxOutConnector[11] = fifoOut[5][8];
              muxOutConnector[12] = fifoOut[6][8];
              muxOutConnector[13] = fifoOut[7][8];
              muxOutConnector[14] = fifoOut[8][8];
              muxOutConnector[15] = fifoOut[9][8];
              muxOutConnector[16] = fifoOut[10][8];
              muxOutConnector[17] = fifoOut[11][8];
              muxOutConnector[18] = fifoOut[12][8];
              muxOutConnector[19] = fifoOut[13][8];
              muxOutConnector[20] = fifoOut[14][8];
              muxOutConnector[21] = fifoOut[15][8];
              muxOutConnector[22] = fifoOut[16][8];
              muxOutConnector[23] = fifoOut[17][8];
              muxOutConnector[24] = fifoOut[18][8];
              muxOutConnector[25] = fifoOut[19][8];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         11: begin
              muxOutConnector[0] = fifoOut[20][9];
              muxOutConnector[1] = fifoOut[21][9];
              muxOutConnector[2] = fifoOut[22][9];
              muxOutConnector[3] = fifoOut[23][9];
              muxOutConnector[4] = fifoOut[24][9];
              muxOutConnector[5] = fifoOut[25][9];
              muxOutConnector[6] = fifoOut[0][8];
              muxOutConnector[7] = fifoOut[1][8];
              muxOutConnector[8] = fifoOut[2][8];
              muxOutConnector[9] = fifoOut[3][8];
              muxOutConnector[10] = fifoOut[4][8];
              muxOutConnector[11] = fifoOut[5][8];
              muxOutConnector[12] = fifoOut[6][8];
              muxOutConnector[13] = fifoOut[7][8];
              muxOutConnector[14] = fifoOut[8][8];
              muxOutConnector[15] = fifoOut[9][8];
              muxOutConnector[16] = fifoOut[10][8];
              muxOutConnector[17] = fifoOut[11][8];
              muxOutConnector[18] = fifoOut[12][8];
              muxOutConnector[19] = fifoOut[13][8];
              muxOutConnector[20] = fifoOut[14][8];
              muxOutConnector[21] = fifoOut[15][8];
              muxOutConnector[22] = fifoOut[16][8];
              muxOutConnector[23] = fifoOut[17][8];
              muxOutConnector[24] = fifoOut[18][8];
              muxOutConnector[25] = fifoOut[19][8];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         12: begin
              muxOutConnector[0] = fifoOut[20][9];
              muxOutConnector[1] = fifoOut[21][9];
              muxOutConnector[2] = fifoOut[22][9];
              muxOutConnector[3] = fifoOut[23][9];
              muxOutConnector[4] = fifoOut[24][9];
              muxOutConnector[5] = fifoOut[25][9];
              muxOutConnector[6] = fifoOut[0][8];
              muxOutConnector[7] = fifoOut[1][8];
              muxOutConnector[8] = fifoOut[2][8];
              muxOutConnector[9] = fifoOut[3][8];
              muxOutConnector[10] = fifoOut[4][8];
              muxOutConnector[11] = fifoOut[5][8];
              muxOutConnector[12] = fifoOut[6][8];
              muxOutConnector[13] = fifoOut[7][8];
              muxOutConnector[14] = fifoOut[8][8];
              muxOutConnector[15] = fifoOut[9][8];
              muxOutConnector[16] = fifoOut[10][8];
              muxOutConnector[17] = fifoOut[11][8];
              muxOutConnector[18] = fifoOut[12][8];
              muxOutConnector[19] = fifoOut[13][8];
              muxOutConnector[20] = fifoOut[14][8];
              muxOutConnector[21] = fifoOut[15][8];
              muxOutConnector[22] = fifoOut[16][8];
              muxOutConnector[23] = fifoOut[17][8];
              muxOutConnector[24] = fifoOut[18][8];
              muxOutConnector[25] = fifoOut[19][8];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         13: begin
              muxOutConnector[0] = fifoOut[20][9];
              muxOutConnector[1] = fifoOut[21][9];
              muxOutConnector[2] = fifoOut[22][9];
              muxOutConnector[3] = fifoOut[23][9];
              muxOutConnector[4] = fifoOut[24][9];
              muxOutConnector[5] = fifoOut[25][9];
              muxOutConnector[6] = fifoOut[0][8];
              muxOutConnector[7] = fifoOut[1][8];
              muxOutConnector[8] = fifoOut[2][8];
              muxOutConnector[9] = fifoOut[3][8];
              muxOutConnector[10] = fifoOut[4][8];
              muxOutConnector[11] = fifoOut[5][8];
              muxOutConnector[12] = fifoOut[6][8];
              muxOutConnector[13] = fifoOut[7][8];
              muxOutConnector[14] = fifoOut[8][8];
              muxOutConnector[15] = fifoOut[9][8];
              muxOutConnector[16] = fifoOut[10][8];
              muxOutConnector[17] = fifoOut[11][8];
              muxOutConnector[18] = fifoOut[12][8];
              muxOutConnector[19] = fifoOut[13][8];
              muxOutConnector[20] = fifoOut[14][8];
              muxOutConnector[21] = fifoOut[15][8];
              muxOutConnector[22] = fifoOut[16][8];
              muxOutConnector[23] = fifoOut[17][8];
              muxOutConnector[24] = fifoOut[18][8];
              muxOutConnector[25] = fifoOut[19][8];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         14: begin
              muxOutConnector[0] = fifoOut[20][9];
              muxOutConnector[1] = fifoOut[21][9];
              muxOutConnector[2] = fifoOut[22][9];
              muxOutConnector[3] = fifoOut[23][9];
              muxOutConnector[4] = fifoOut[24][9];
              muxOutConnector[5] = fifoOut[25][9];
              muxOutConnector[6] = fifoOut[0][8];
              muxOutConnector[7] = fifoOut[1][8];
              muxOutConnector[8] = fifoOut[26][12];
              muxOutConnector[9] = fifoOut[27][12];
              muxOutConnector[10] = fifoOut[28][12];
              muxOutConnector[11] = fifoOut[29][12];
              muxOutConnector[12] = fifoOut[30][12];
              muxOutConnector[13] = fifoOut[31][12];
              muxOutConnector[14] = fifoOut[32][12];
              muxOutConnector[15] = fifoOut[33][12];
              muxOutConnector[16] = fifoOut[34][12];
              muxOutConnector[17] = fifoOut[35][12];
              muxOutConnector[18] = fifoOut[36][12];
              muxOutConnector[19] = fifoOut[37][12];
              muxOutConnector[20] = fifoOut[38][12];
              muxOutConnector[21] = fifoOut[39][12];
              muxOutConnector[22] = fifoOut[40][12];
              muxOutConnector[23] = fifoOut[41][12];
              muxOutConnector[24] = fifoOut[42][12];
              muxOutConnector[25] = fifoOut[43][12];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         15: begin
              muxOutConnector[0] = fifoOut[44][13];
              muxOutConnector[1] = fifoOut[45][13];
              muxOutConnector[2] = fifoOut[46][13];
              muxOutConnector[3] = fifoOut[47][13];
              muxOutConnector[4] = fifoOut[48][13];
              muxOutConnector[5] = fifoOut[49][13];
              muxOutConnector[6] = fifoOut[50][13];
              muxOutConnector[7] = fifoOut[51][13];
              muxOutConnector[8] = fifoOut[26][12];
              muxOutConnector[9] = fifoOut[27][12];
              muxOutConnector[10] = fifoOut[28][12];
              muxOutConnector[11] = fifoOut[29][12];
              muxOutConnector[12] = fifoOut[30][12];
              muxOutConnector[13] = fifoOut[31][12];
              muxOutConnector[14] = fifoOut[32][12];
              muxOutConnector[15] = fifoOut[33][12];
              muxOutConnector[16] = fifoOut[34][12];
              muxOutConnector[17] = fifoOut[35][12];
              muxOutConnector[18] = fifoOut[36][12];
              muxOutConnector[19] = fifoOut[37][12];
              muxOutConnector[20] = fifoOut[38][12];
              muxOutConnector[21] = fifoOut[39][12];
              muxOutConnector[22] = fifoOut[40][12];
              muxOutConnector[23] = fifoOut[41][12];
              muxOutConnector[24] = fifoOut[42][12];
              muxOutConnector[25] = fifoOut[43][12];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[17][16];
              muxOutConnector[29] = fifoOut[18][16];
              muxOutConnector[30] = fifoOut[19][16];
              muxOutConnector[31] = fifoOut[20][16];
              muxOutConnector[32] = fifoOut[21][16];
              muxOutConnector[33] = fifoOut[22][16];
              muxOutConnector[34] = fifoOut[23][16];
              muxOutConnector[35] = fifoOut[24][16];
              muxOutConnector[36] = fifoOut[25][16];
              muxOutConnector[37] = fifoOut[0][15];
              muxOutConnector[38] = fifoOut[1][15];
              muxOutConnector[39] = fifoOut[2][15];
              muxOutConnector[40] = fifoOut[3][15];
              muxOutConnector[41] = fifoOut[4][15];
              muxOutConnector[42] = fifoOut[5][15];
              muxOutConnector[43] = fifoOut[6][15];
              muxOutConnector[44] = fifoOut[7][15];
              muxOutConnector[45] = fifoOut[8][15];
              muxOutConnector[46] = fifoOut[9][15];
              muxOutConnector[47] = fifoOut[10][15];
              muxOutConnector[48] = fifoOut[11][15];
              muxOutConnector[49] = fifoOut[12][15];
              muxOutConnector[50] = fifoOut[13][15];
              muxOutConnector[51] = fifoOut[14][15];
         end
         16: begin
              muxOutConnector[0] = fifoOut[44][13];
              muxOutConnector[1] = fifoOut[45][13];
              muxOutConnector[2] = fifoOut[46][13];
              muxOutConnector[3] = fifoOut[47][13];
              muxOutConnector[4] = fifoOut[48][13];
              muxOutConnector[5] = fifoOut[49][13];
              muxOutConnector[6] = fifoOut[50][13];
              muxOutConnector[7] = fifoOut[51][13];
              muxOutConnector[8] = fifoOut[26][12];
              muxOutConnector[9] = fifoOut[27][12];
              muxOutConnector[10] = fifoOut[28][12];
              muxOutConnector[11] = fifoOut[29][12];
              muxOutConnector[12] = fifoOut[30][12];
              muxOutConnector[13] = fifoOut[31][12];
              muxOutConnector[14] = fifoOut[32][12];
              muxOutConnector[15] = fifoOut[33][12];
              muxOutConnector[16] = fifoOut[34][12];
              muxOutConnector[17] = fifoOut[35][12];
              muxOutConnector[18] = fifoOut[36][12];
              muxOutConnector[19] = fifoOut[37][12];
              muxOutConnector[20] = fifoOut[38][12];
              muxOutConnector[21] = fifoOut[39][12];
              muxOutConnector[22] = fifoOut[40][12];
              muxOutConnector[23] = fifoOut[41][12];
              muxOutConnector[24] = fifoOut[42][12];
              muxOutConnector[25] = fifoOut[43][12];
              muxOutConnector[26] = fifoOut[15][16];
              muxOutConnector[27] = fifoOut[16][16];
              muxOutConnector[28] = fifoOut[41][3];
              muxOutConnector[29] = fifoOut[42][3];
              muxOutConnector[30] = fifoOut[43][3];
              muxOutConnector[31] = fifoOut[44][3];
              muxOutConnector[32] = fifoOut[45][3];
              muxOutConnector[33] = fifoOut[46][3];
              muxOutConnector[34] = fifoOut[47][3];
              muxOutConnector[35] = fifoOut[48][3];
              muxOutConnector[36] = fifoOut[49][3];
              muxOutConnector[37] = fifoOut[50][3];
              muxOutConnector[38] = fifoOut[51][3];
              muxOutConnector[39] = fifoOut[26][2];
              muxOutConnector[40] = fifoOut[27][2];
              muxOutConnector[41] = fifoOut[28][2];
              muxOutConnector[42] = fifoOut[29][2];
              muxOutConnector[43] = fifoOut[30][2];
              muxOutConnector[44] = fifoOut[31][2];
              muxOutConnector[45] = fifoOut[32][2];
              muxOutConnector[46] = fifoOut[33][2];
              muxOutConnector[47] = fifoOut[34][2];
              muxOutConnector[48] = fifoOut[35][2];
              muxOutConnector[49] = fifoOut[36][2];
              muxOutConnector[50] = fifoOut[37][2];
              muxOutConnector[51] = fifoOut[38][2];
         end
         17: begin
              muxOutConnector[0] = fifoOut[44][13];
              muxOutConnector[1] = fifoOut[45][13];
              muxOutConnector[2] = fifoOut[46][13];
              muxOutConnector[3] = fifoOut[47][13];
              muxOutConnector[4] = fifoOut[48][13];
              muxOutConnector[5] = fifoOut[49][13];
              muxOutConnector[6] = fifoOut[50][13];
              muxOutConnector[7] = fifoOut[51][13];
              muxOutConnector[8] = fifoOut[26][12];
              muxOutConnector[9] = fifoOut[27][12];
              muxOutConnector[10] = fifoOut[28][12];
              muxOutConnector[11] = fifoOut[29][12];
              muxOutConnector[12] = fifoOut[30][12];
              muxOutConnector[13] = fifoOut[31][12];
              muxOutConnector[14] = fifoOut[32][12];
              muxOutConnector[15] = fifoOut[33][12];
              muxOutConnector[16] = fifoOut[34][12];
              muxOutConnector[17] = fifoOut[35][12];
              muxOutConnector[18] = fifoOut[36][12];
              muxOutConnector[19] = fifoOut[37][12];
              muxOutConnector[20] = fifoOut[38][12];
              muxOutConnector[21] = fifoOut[39][12];
              muxOutConnector[22] = fifoOut[40][12];
              muxOutConnector[23] = fifoOut[41][12];
              muxOutConnector[24] = fifoOut[42][12];
              muxOutConnector[25] = fifoOut[43][12];
              muxOutConnector[26] = fifoOut[39][3];
              muxOutConnector[27] = fifoOut[40][3];
              muxOutConnector[28] = fifoOut[41][3];
              muxOutConnector[29] = fifoOut[42][3];
              muxOutConnector[30] = fifoOut[43][3];
              muxOutConnector[31] = fifoOut[44][3];
              muxOutConnector[32] = fifoOut[45][3];
              muxOutConnector[33] = fifoOut[46][3];
              muxOutConnector[34] = fifoOut[47][3];
              muxOutConnector[35] = fifoOut[48][3];
              muxOutConnector[36] = fifoOut[49][3];
              muxOutConnector[37] = fifoOut[50][3];
              muxOutConnector[38] = fifoOut[51][3];
              muxOutConnector[39] = fifoOut[26][2];
              muxOutConnector[40] = fifoOut[27][2];
              muxOutConnector[41] = fifoOut[28][2];
              muxOutConnector[42] = fifoOut[29][2];
              muxOutConnector[43] = fifoOut[30][2];
              muxOutConnector[44] = fifoOut[31][2];
              muxOutConnector[45] = fifoOut[32][2];
              muxOutConnector[46] = fifoOut[33][2];
              muxOutConnector[47] = fifoOut[34][2];
              muxOutConnector[48] = fifoOut[35][2];
              muxOutConnector[49] = fifoOut[36][2];
              muxOutConnector[50] = fifoOut[37][2];
              muxOutConnector[51] = fifoOut[38][2];
         end
         18: begin
              muxOutConnector[0] = fifoOut[44][13];
              muxOutConnector[1] = fifoOut[45][13];
              muxOutConnector[2] = fifoOut[46][13];
              muxOutConnector[3] = fifoOut[47][13];
              muxOutConnector[4] = fifoOut[48][13];
              muxOutConnector[5] = fifoOut[49][13];
              muxOutConnector[6] = fifoOut[50][13];
              muxOutConnector[7] = fifoOut[51][13];
              muxOutConnector[8] = fifoOut[26][12];
              muxOutConnector[9] = fifoOut[27][12];
              muxOutConnector[10] = fifoOut[28][12];
              muxOutConnector[11] = fifoOut[29][12];
              muxOutConnector[12] = fifoOut[30][12];
              muxOutConnector[13] = fifoOut[31][12];
              muxOutConnector[14] = fifoOut[32][12];
              muxOutConnector[15] = fifoOut[33][12];
              muxOutConnector[16] = fifoOut[34][12];
              muxOutConnector[17] = fifoOut[35][12];
              muxOutConnector[18] = fifoOut[36][12];
              muxOutConnector[19] = fifoOut[37][12];
              muxOutConnector[20] = fifoOut[38][12];
              muxOutConnector[21] = fifoOut[39][12];
              muxOutConnector[22] = fifoOut[40][12];
              muxOutConnector[23] = fifoOut[41][12];
              muxOutConnector[24] = fifoOut[42][12];
              muxOutConnector[25] = fifoOut[43][12];
              muxOutConnector[26] = fifoOut[39][3];
              muxOutConnector[27] = fifoOut[40][3];
              muxOutConnector[28] = fifoOut[41][3];
              muxOutConnector[29] = fifoOut[42][3];
              muxOutConnector[30] = fifoOut[43][3];
              muxOutConnector[31] = fifoOut[44][3];
              muxOutConnector[32] = fifoOut[45][3];
              muxOutConnector[33] = fifoOut[46][3];
              muxOutConnector[34] = fifoOut[47][3];
              muxOutConnector[35] = fifoOut[48][3];
              muxOutConnector[36] = fifoOut[49][3];
              muxOutConnector[37] = fifoOut[50][3];
              muxOutConnector[38] = fifoOut[51][3];
              muxOutConnector[39] = fifoOut[26][2];
              muxOutConnector[40] = fifoOut[27][2];
              muxOutConnector[41] = fifoOut[28][2];
              muxOutConnector[42] = fifoOut[29][2];
              muxOutConnector[43] = fifoOut[30][2];
              muxOutConnector[44] = fifoOut[31][2];
              muxOutConnector[45] = fifoOut[32][2];
              muxOutConnector[46] = fifoOut[33][2];
              muxOutConnector[47] = fifoOut[34][2];
              muxOutConnector[48] = fifoOut[35][2];
              muxOutConnector[49] = fifoOut[36][2];
              muxOutConnector[50] = fifoOut[37][2];
              muxOutConnector[51] = fifoOut[38][2];
         end
         19: begin
              muxOutConnector[0] = fifoOut[44][13];
              muxOutConnector[1] = fifoOut[45][13];
              muxOutConnector[2] = fifoOut[46][13];
              muxOutConnector[3] = fifoOut[47][13];
              muxOutConnector[4] = fifoOut[48][13];
              muxOutConnector[5] = fifoOut[49][13];
              muxOutConnector[6] = fifoOut[50][13];
              muxOutConnector[7] = fifoOut[51][13];
              muxOutConnector[8] = fifoOut[26][12];
              muxOutConnector[9] = fifoOut[27][12];
              muxOutConnector[10] = fifoOut[28][12];
              muxOutConnector[11] = fifoOut[29][12];
              muxOutConnector[12] = fifoOut[30][12];
              muxOutConnector[13] = fifoOut[31][12];
              muxOutConnector[14] = fifoOut[32][12];
              muxOutConnector[15] = fifoOut[33][12];
              muxOutConnector[16] = fifoOut[34][12];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[39][3];
              muxOutConnector[27] = fifoOut[40][3];
              muxOutConnector[28] = fifoOut[41][3];
              muxOutConnector[29] = fifoOut[42][3];
              muxOutConnector[30] = fifoOut[43][3];
              muxOutConnector[31] = fifoOut[44][3];
              muxOutConnector[32] = fifoOut[45][3];
              muxOutConnector[33] = fifoOut[46][3];
              muxOutConnector[34] = fifoOut[47][3];
              muxOutConnector[35] = fifoOut[48][3];
              muxOutConnector[36] = fifoOut[49][3];
              muxOutConnector[37] = fifoOut[50][3];
              muxOutConnector[38] = fifoOut[51][3];
              muxOutConnector[39] = fifoOut[26][2];
              muxOutConnector[40] = fifoOut[27][2];
              muxOutConnector[41] = fifoOut[28][2];
              muxOutConnector[42] = fifoOut[29][2];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
         end
         default: begin
               for(i=0;i<muxOutSymbols;i=i+1)begin
                muxOutConnector[i] = 0;
              end
         end
//hgjhgbuiguigbigbgbgbui
         endcase
    end
endcase
             end
        endmodule