`timescale 1ns / 1ps
module Dmem_circ9_scripted(
		 muxOut,
		 dMemIn,
		 wr_en,
		 reaccessAddress,
		 reaccess_lyr,
		 rd_en, clk, rst 
 );
parameter r = 52;
parameter c = 12;
parameter w = 6;
parameter ADDRESSWIDTH = 5;

parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 
output wire [r*w -1 : 0]muxOut;// r numbers of w bits
input [r*w-1:0]dMemIn;
input wr_en;
input [ADDRESSWIDTH-1:0]reaccessAddress;
input reaccess_lyr;
input rd_en;
input clk,rst;

wire [(ADDRESSWIDTH+1)-1:0]case_sel;//{layer,address}
wire [w-1:0]dMemInDummy[r-1:0];
reg [w-1:0]muxOutWire[r-1:0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<r;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutWire[k];
        assign dMemInDummy[k] = dMemIn[ (k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always @(posedge clk) begin
    if (rst) begin
         for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] = 0;
           end
        end
    end
    else begin
    if(wr_en) begin
        // Set (i,j)th value = (i,j-1)th value
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Load Inputs
        for(i = r-1; i > -1; i=i-1) begin
            fifoOut[i][0] <= dMemInDummy[i]; 
        end
    end
    else begin 
        // Set (i,j)th value = (i,j)th value
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <= fifoOut[i][j];
            end
        end
    end
    end
end

assign case_sel = rd_en ? {reaccess_lyr,reaccessAddress} : {1'd1,READDISABLEDCASE};

always@(*) begin
    case(case_sel)

		 {1'd0, 5'd0} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd1} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd2} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd3} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd4} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd5} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd6} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd7} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd8} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd9} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 3 ][ 6 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 4 ][ 6 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 5 ][ 6 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 6 ][ 6 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 7 ][ 6 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 8 ][ 6 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 9 ][ 6 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 10 ][ 6 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 11 ][ 6 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 12 ][ 6 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 13 ][ 6 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 14 ][ 6 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 15 ][ 6 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 16 ][ 6 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 17 ][ 6 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 18 ][ 6 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 19 ][ 6 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 20 ][ 6 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 21 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 22 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 23 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 24 ][ 6 ]; 
		 end
		 {1'd0, 5'd10} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = fifoOut[ 26 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 27 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 28 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 29 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 30 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 3 ][ 6 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 4 ][ 6 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 5 ][ 6 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 6 ][ 6 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 7 ][ 6 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 8 ][ 6 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 9 ][ 6 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 10 ][ 6 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 11 ][ 6 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 12 ][ 6 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 13 ][ 6 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 14 ][ 6 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 15 ][ 6 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 16 ][ 6 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 17 ][ 6 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 18 ][ 6 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 19 ][ 6 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 20 ][ 6 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 21 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 22 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 23 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 24 ][ 6 ]; 
		 end
		 {1'd0, 5'd11} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 36 ][ 8 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 37 ][ 8 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 38 ][ 8 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 39 ][ 8 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 40 ][ 8 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 41 ][ 8 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 42 ][ 8 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 43 ][ 8 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 44 ][ 8 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 45 ][ 8 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 46 ][ 8 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 47 ][ 8 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 48 ][ 8 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 49 ][ 8 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 50 ][ 8 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 51 ][ 8 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 26 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 27 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 28 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 29 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 30 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 3 ][ 6 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 4 ][ 6 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 5 ][ 6 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 6 ][ 6 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 7 ][ 6 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 8 ][ 6 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 9 ][ 6 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 10 ][ 6 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 11 ][ 6 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 12 ][ 6 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 13 ][ 6 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 14 ][ 6 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 15 ][ 6 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 16 ][ 6 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 17 ][ 6 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 18 ][ 6 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 19 ][ 6 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 20 ][ 6 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 21 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 22 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 23 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 24 ][ 6 ]; 
		 end
		 {1'd0, 5'd12} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 36 ][ 8 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 37 ][ 8 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 38 ][ 8 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 39 ][ 8 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 40 ][ 8 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 41 ][ 8 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 42 ][ 8 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 43 ][ 8 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 44 ][ 8 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 45 ][ 8 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 46 ][ 8 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 47 ][ 8 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 48 ][ 8 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 49 ][ 8 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 50 ][ 8 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 51 ][ 8 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 26 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 27 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 28 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 29 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 30 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 3 ][ 6 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 4 ][ 6 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 5 ][ 6 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 6 ][ 6 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 7 ][ 6 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 8 ][ 6 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 9 ][ 6 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 10 ][ 6 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 11 ][ 6 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 12 ][ 6 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 13 ][ 6 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 14 ][ 6 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 15 ][ 6 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 16 ][ 6 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 17 ][ 6 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 18 ][ 6 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 19 ][ 6 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 20 ][ 6 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 21 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 22 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 23 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 24 ][ 6 ]; 
		 end
		 {1'd0, 5'd13} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 36 ][ 8 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 37 ][ 8 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 38 ][ 8 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 39 ][ 8 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 40 ][ 8 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 41 ][ 8 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 42 ][ 8 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 43 ][ 8 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 44 ][ 8 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 45 ][ 8 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 46 ][ 8 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 47 ][ 8 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 48 ][ 8 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 49 ][ 8 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 50 ][ 8 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 51 ][ 8 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 26 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 27 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 28 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 29 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 30 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 3 ][ 6 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 4 ][ 6 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 5 ][ 6 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 6 ][ 6 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 7 ][ 6 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 8 ][ 6 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 9 ][ 6 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 10 ][ 6 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 11 ][ 6 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 12 ][ 6 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 13 ][ 6 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 14 ][ 6 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 15 ][ 6 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 16 ][ 6 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 17 ][ 6 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 18 ][ 6 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 19 ][ 6 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 20 ][ 6 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 21 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 22 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 23 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 24 ][ 6 ]; 
		 end
		 {1'd0, 5'd14} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 36 ][ 8 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 37 ][ 8 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 38 ][ 8 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 39 ][ 8 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 40 ][ 8 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 41 ][ 8 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 42 ][ 8 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 43 ][ 8 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 44 ][ 8 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 45 ][ 8 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 46 ][ 8 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 47 ][ 8 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 48 ][ 8 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 49 ][ 8 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 50 ][ 8 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 51 ][ 8 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 26 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 27 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 28 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 29 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 30 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 3 ][ 6 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 4 ][ 6 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 5 ][ 6 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 6 ][ 6 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 7 ][ 6 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 8 ][ 6 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 9 ][ 6 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 10 ][ 6 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 11 ][ 6 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 12 ][ 6 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 13 ][ 6 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 14 ][ 6 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 15 ][ 6 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 16 ][ 6 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 17 ][ 6 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 18 ][ 6 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 19 ][ 6 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 20 ][ 6 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 21 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 22 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 23 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 24 ][ 6 ]; 
		 end
		 {1'd0, 5'd15} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 36 ][ 8 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 37 ][ 8 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 38 ][ 8 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 39 ][ 8 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 40 ][ 8 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 41 ][ 8 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 42 ][ 8 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 43 ][ 8 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 44 ][ 8 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 45 ][ 8 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 46 ][ 8 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 47 ][ 8 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 48 ][ 8 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 49 ][ 8 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 50 ][ 8 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 51 ][ 8 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 26 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 27 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 28 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 29 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 30 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 3 ][ 6 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 4 ][ 6 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 5 ][ 6 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 6 ][ 6 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 7 ][ 6 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 8 ][ 6 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 9 ][ 6 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 10 ][ 6 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 11 ][ 6 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 12 ][ 6 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 13 ][ 6 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 14 ][ 6 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 15 ][ 6 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 16 ][ 6 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 17 ][ 6 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 18 ][ 6 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 19 ][ 6 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 20 ][ 6 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 21 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 22 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 23 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 24 ][ 6 ]; 
		 end
		 {1'd0, 5'd16} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 36 ][ 8 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 37 ][ 8 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 38 ][ 8 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 39 ][ 8 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 40 ][ 8 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 41 ][ 8 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 42 ][ 8 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 43 ][ 8 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 44 ][ 8 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 45 ][ 8 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 46 ][ 8 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 47 ][ 8 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 48 ][ 8 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 49 ][ 8 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 50 ][ 8 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 51 ][ 8 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 26 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 27 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 28 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 29 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 30 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 3 ][ 6 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 4 ][ 6 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 5 ][ 6 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 6 ][ 6 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 7 ][ 6 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 8 ][ 6 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 9 ][ 6 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 10 ][ 6 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 11 ][ 6 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 12 ][ 6 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 13 ][ 6 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 14 ][ 6 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 15 ][ 6 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 16 ][ 6 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 17 ][ 6 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 18 ][ 6 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 19 ][ 6 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 20 ][ 6 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 21 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 22 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 23 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 24 ][ 6 ]; 
		 end
		 {1'd0, 5'd17} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 36 ][ 8 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 37 ][ 8 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 38 ][ 8 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 39 ][ 8 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 40 ][ 8 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 41 ][ 8 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 42 ][ 8 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 43 ][ 8 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 44 ][ 8 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 45 ][ 8 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 46 ][ 8 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 47 ][ 8 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 48 ][ 8 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 49 ][ 8 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 50 ][ 8 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 51 ][ 8 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 26 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 27 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 28 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 29 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 30 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 3 ][ 6 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 4 ][ 6 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 5 ][ 6 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 6 ][ 6 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 7 ][ 6 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 8 ][ 6 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 9 ][ 6 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 10 ][ 6 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 11 ][ 6 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 12 ][ 6 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 13 ][ 6 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 14 ][ 6 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 15 ][ 6 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 16 ][ 6 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 17 ][ 6 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 18 ][ 6 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 19 ][ 6 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 20 ][ 6 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 21 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 22 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 23 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 24 ][ 6 ]; 
		 end
		 {1'd0, 5'd18} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 36 ][ 8 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 37 ][ 8 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 38 ][ 8 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 39 ][ 8 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 40 ][ 8 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 41 ][ 8 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 42 ][ 8 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 43 ][ 8 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 44 ][ 8 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 45 ][ 8 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 46 ][ 8 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 47 ][ 8 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 48 ][ 8 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 49 ][ 8 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 50 ][ 8 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 51 ][ 8 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 26 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 27 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 28 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 29 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 30 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 3 ][ 6 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 4 ][ 6 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 5 ][ 6 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 6 ][ 6 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 7 ][ 6 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 8 ][ 6 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 9 ][ 6 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 10 ][ 6 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 11 ][ 6 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 12 ][ 6 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 13 ][ 6 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 14 ][ 6 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 15 ][ 6 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 16 ][ 6 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 17 ][ 6 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 18 ][ 6 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 19 ][ 6 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 20 ][ 6 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 21 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 22 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 23 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 24 ][ 6 ]; 
		 end
		 {1'd0, 5'd19} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 36 ][ 8 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 37 ][ 8 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 38 ][ 8 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 39 ][ 8 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 40 ][ 8 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 41 ][ 8 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 42 ][ 8 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 43 ][ 8 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 44 ][ 8 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 45 ][ 8 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 46 ][ 8 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 47 ][ 8 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 48 ][ 8 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 49 ][ 8 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 50 ][ 8 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 51 ][ 8 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 26 ][ 7 ]; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 3 ][ 6 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 4 ][ 6 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 5 ][ 6 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 6 ][ 6 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 7 ][ 6 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 8 ][ 6 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 9 ][ 6 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 10 ][ 6 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 11 ][ 6 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 12 ][ 6 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 13 ][ 6 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 14 ][ 6 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 15 ][ 6 ]; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd0} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd1} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd2} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd3} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd4} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd5} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = fifoOut[ 26 ][ 2 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 27 ][ 2 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 28 ][ 2 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 29 ][ 2 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 30 ][ 2 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 31 ][ 2 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 32 ][ 2 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd6} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 51 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 26 ][ 2 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 27 ][ 2 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 28 ][ 2 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 29 ][ 2 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 30 ][ 2 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 31 ][ 2 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 32 ][ 2 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd7} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 51 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 26 ][ 2 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 27 ][ 2 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 28 ][ 2 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 29 ][ 2 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 30 ][ 2 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 31 ][ 2 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 32 ][ 2 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd8} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 51 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 26 ][ 2 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 27 ][ 2 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 28 ][ 2 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 29 ][ 2 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 30 ][ 2 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 31 ][ 2 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 32 ][ 2 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd9} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 51 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 26 ][ 2 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 27 ][ 2 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 28 ][ 2 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 29 ][ 2 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 30 ][ 2 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 31 ][ 2 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 32 ][ 2 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd10} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 51 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 26 ][ 2 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 27 ][ 2 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 28 ][ 2 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 29 ][ 2 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 30 ][ 2 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 31 ][ 2 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 32 ][ 2 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd11} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 51 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 26 ][ 2 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 27 ][ 2 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 28 ][ 2 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 29 ][ 2 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 30 ][ 2 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 31 ][ 2 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 32 ][ 2 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd12} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 51 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 26 ][ 2 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 27 ][ 2 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 28 ][ 2 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 29 ][ 2 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 30 ][ 2 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 31 ][ 2 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 32 ][ 2 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd13} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 51 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 26 ][ 2 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 27 ][ 2 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 28 ][ 2 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 29 ][ 2 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 30 ][ 2 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 31 ][ 2 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 32 ][ 2 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = fifoOut[ 0 ][ 10 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 1 ][ 10 ]; 
		 end
		 {1'd1, 5'd14} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 51 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 26 ][ 2 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 27 ][ 2 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 28 ][ 2 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 29 ][ 2 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 30 ][ 2 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 31 ][ 2 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 32 ][ 2 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 2 ][ 11 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 3 ][ 11 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 4 ][ 11 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 5 ][ 11 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 6 ][ 11 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 7 ][ 11 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 8 ][ 11 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 9 ][ 11 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 10 ][ 11 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 11 ][ 11 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 12 ][ 11 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 13 ][ 11 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 14 ][ 11 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 15 ][ 11 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 16 ][ 11 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 17 ][ 11 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 18 ][ 11 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 19 ][ 11 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 20 ][ 11 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 21 ][ 11 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 22 ][ 11 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 23 ][ 11 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 24 ][ 11 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 25 ][ 11 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 0 ][ 10 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 1 ][ 10 ]; 
		 end
		 {1'd1, 5'd15} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 51 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 26 ][ 2 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 27 ][ 2 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 28 ][ 2 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 29 ][ 2 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 30 ][ 2 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 31 ][ 2 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 32 ][ 2 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 2 ][ 11 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 3 ][ 11 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 4 ][ 11 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 5 ][ 11 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 6 ][ 11 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 7 ][ 11 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 8 ][ 11 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 9 ][ 11 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 10 ][ 11 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 11 ][ 11 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 12 ][ 11 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 13 ][ 11 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 14 ][ 11 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 15 ][ 11 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 16 ][ 11 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 17 ][ 11 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 18 ][ 11 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 19 ][ 11 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 20 ][ 11 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 21 ][ 11 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 22 ][ 11 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 23 ][ 11 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 24 ][ 11 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 25 ][ 11 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 0 ][ 10 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 1 ][ 10 ]; 
		 end
		 {1'd1, 5'd16} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 51 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 26 ][ 2 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 27 ][ 2 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 28 ][ 2 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 29 ][ 2 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 30 ][ 2 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 31 ][ 2 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 32 ][ 2 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 2 ][ 11 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 3 ][ 11 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 4 ][ 11 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 5 ][ 11 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 6 ][ 11 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 7 ][ 11 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 8 ][ 11 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 9 ][ 11 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 10 ][ 11 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 11 ][ 11 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 12 ][ 11 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 13 ][ 11 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 14 ][ 11 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 15 ][ 11 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 16 ][ 11 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 17 ][ 11 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 18 ][ 11 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 19 ][ 11 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 20 ][ 11 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 21 ][ 11 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 22 ][ 11 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 23 ][ 11 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 24 ][ 11 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 25 ][ 11 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 0 ][ 10 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 1 ][ 10 ]; 
		 end
		 {1'd1, 5'd17} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 51 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 26 ][ 2 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 27 ][ 2 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 28 ][ 2 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 29 ][ 2 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 30 ][ 2 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 31 ][ 2 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 32 ][ 2 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 2 ][ 11 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 3 ][ 11 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 4 ][ 11 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 5 ][ 11 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 6 ][ 11 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 7 ][ 11 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 8 ][ 11 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 9 ][ 11 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 10 ][ 11 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 11 ][ 11 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 12 ][ 11 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 13 ][ 11 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 14 ][ 11 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 15 ][ 11 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 16 ][ 11 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 17 ][ 11 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 18 ][ 11 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 19 ][ 11 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 20 ][ 11 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 21 ][ 11 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 22 ][ 11 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 23 ][ 11 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 24 ][ 11 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 25 ][ 11 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 0 ][ 10 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 1 ][ 10 ]; 
		 end
		 {1'd1, 5'd18} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 51 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 26 ][ 2 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 27 ][ 2 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 28 ][ 2 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 29 ][ 2 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 30 ][ 2 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 31 ][ 2 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 32 ][ 2 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 2 ][ 11 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 3 ][ 11 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 4 ][ 11 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 5 ][ 11 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 6 ][ 11 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 7 ][ 11 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 8 ][ 11 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 9 ][ 11 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 10 ][ 11 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 11 ][ 11 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 12 ][ 11 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 13 ][ 11 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 14 ][ 11 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 15 ][ 11 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 16 ][ 11 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 17 ][ 11 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 18 ][ 11 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 19 ][ 11 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 20 ][ 11 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 21 ][ 11 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 22 ][ 11 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 23 ][ 11 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 24 ][ 11 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 25 ][ 11 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 0 ][ 10 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 1 ][ 10 ]; 
		 end
		 {1'd1, 5'd19} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 2 ][ 11 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 3 ][ 11 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 4 ][ 11 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 5 ][ 11 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 6 ][ 11 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 7 ][ 11 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 8 ][ 11 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 9 ][ 11 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 10 ][ 11 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 11 ][ 11 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 12 ][ 11 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 13 ][ 11 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 14 ][ 11 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 15 ][ 11 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 16 ][ 11 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 17 ][ 11 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 18 ][ 11 ]; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
    default:begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
    end
    endcase
end
endmodule
