`timescale 1ns / 1ps
module LMem1To0_511_circ11_ys_yu_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        wr_en,
        feedback_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 13;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input [ADDRESSWIDTH-1:0]unloadAddress;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

input feedback_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        if(feedback_en) begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= fifoOut[i][c-1];
         end
        end
        else begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= ly0InConnector[i];
         end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
       0: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = fifoOut[8][7][w-1];
              unloadMuxOut[22] = fifoOut[9][7][w-1];
              unloadMuxOut[23] = fifoOut[10][7][w-1];
              unloadMuxOut[24] = fifoOut[11][7][w-1];
              unloadMuxOut[25] = fifoOut[12][7][w-1];
              unloadMuxOut[26] = fifoOut[13][7][w-1];
              unloadMuxOut[27] = fifoOut[14][7][w-1];
              unloadMuxOut[28] = fifoOut[15][7][w-1];
              unloadMuxOut[29] = fifoOut[16][7][w-1];
              unloadMuxOut[30] = fifoOut[17][7][w-1];
              unloadMuxOut[31] = fifoOut[18][7][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[19][7][w-1];
              unloadMuxOut[1] = fifoOut[20][7][w-1];
              unloadMuxOut[2] = fifoOut[21][7][w-1];
              unloadMuxOut[3] = fifoOut[22][7][w-1];
              unloadMuxOut[4] = fifoOut[23][7][w-1];
              unloadMuxOut[5] = fifoOut[24][7][w-1];
              unloadMuxOut[6] = fifoOut[25][7][w-1];
              unloadMuxOut[7] = fifoOut[0][6][w-1];
              unloadMuxOut[8] = fifoOut[1][6][w-1];
              unloadMuxOut[9] = fifoOut[2][6][w-1];
              unloadMuxOut[10] = fifoOut[3][6][w-1];
              unloadMuxOut[11] = fifoOut[4][6][w-1];
              unloadMuxOut[12] = fifoOut[5][6][w-1];
              unloadMuxOut[13] = fifoOut[6][6][w-1];
              unloadMuxOut[14] = fifoOut[7][6][w-1];
              unloadMuxOut[15] = fifoOut[8][6][w-1];
              unloadMuxOut[16] = fifoOut[9][6][w-1];
              unloadMuxOut[17] = fifoOut[10][6][w-1];
              unloadMuxOut[18] = fifoOut[11][6][w-1];
              unloadMuxOut[19] = fifoOut[12][6][w-1];
              unloadMuxOut[20] = fifoOut[13][6][w-1];
              unloadMuxOut[21] = fifoOut[14][6][w-1];
              unloadMuxOut[22] = fifoOut[15][6][w-1];
              unloadMuxOut[23] = fifoOut[16][6][w-1];
              unloadMuxOut[24] = fifoOut[17][6][w-1];
              unloadMuxOut[25] = fifoOut[18][6][w-1];
              unloadMuxOut[26] = fifoOut[19][6][w-1];
              unloadMuxOut[27] = fifoOut[20][6][w-1];
              unloadMuxOut[28] = fifoOut[21][6][w-1];
              unloadMuxOut[29] = fifoOut[22][6][w-1];
              unloadMuxOut[30] = fifoOut[23][6][w-1];
              unloadMuxOut[31] = fifoOut[24][6][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[25][6][w-1];
              unloadMuxOut[1] = fifoOut[0][5][w-1];
              unloadMuxOut[2] = fifoOut[1][5][w-1];
              unloadMuxOut[3] = fifoOut[2][5][w-1];
              unloadMuxOut[4] = fifoOut[3][5][w-1];
              unloadMuxOut[5] = fifoOut[4][5][w-1];
              unloadMuxOut[6] = fifoOut[5][5][w-1];
              unloadMuxOut[7] = fifoOut[6][5][w-1];
              unloadMuxOut[8] = fifoOut[7][5][w-1];
              unloadMuxOut[9] = fifoOut[8][5][w-1];
              unloadMuxOut[10] = fifoOut[9][5][w-1];
              unloadMuxOut[11] = fifoOut[10][5][w-1];
              unloadMuxOut[12] = fifoOut[11][5][w-1];
              unloadMuxOut[13] = fifoOut[12][5][w-1];
              unloadMuxOut[14] = fifoOut[26][12][w-1];
              unloadMuxOut[15] = fifoOut[27][12][w-1];
              unloadMuxOut[16] = fifoOut[28][12][w-1];
              unloadMuxOut[17] = fifoOut[29][12][w-1];
              unloadMuxOut[18] = fifoOut[30][12][w-1];
              unloadMuxOut[19] = fifoOut[31][12][w-1];
              unloadMuxOut[20] = fifoOut[32][12][w-1];
              unloadMuxOut[21] = fifoOut[33][12][w-1];
              unloadMuxOut[22] = fifoOut[34][12][w-1];
              unloadMuxOut[23] = fifoOut[35][12][w-1];
              unloadMuxOut[24] = fifoOut[36][12][w-1];
              unloadMuxOut[25] = fifoOut[37][12][w-1];
              unloadMuxOut[26] = fifoOut[38][12][w-1];
              unloadMuxOut[27] = fifoOut[39][12][w-1];
              unloadMuxOut[28] = fifoOut[40][12][w-1];
              unloadMuxOut[29] = fifoOut[41][12][w-1];
              unloadMuxOut[30] = fifoOut[42][12][w-1];
              unloadMuxOut[31] = fifoOut[43][12][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[44][12][w-1];
              unloadMuxOut[1] = fifoOut[45][12][w-1];
              unloadMuxOut[2] = fifoOut[46][12][w-1];
              unloadMuxOut[3] = fifoOut[47][12][w-1];
              unloadMuxOut[4] = fifoOut[48][12][w-1];
              unloadMuxOut[5] = fifoOut[49][12][w-1];
              unloadMuxOut[6] = fifoOut[50][12][w-1];
              unloadMuxOut[7] = fifoOut[51][12][w-1];
              unloadMuxOut[8] = fifoOut[26][11][w-1];
              unloadMuxOut[9] = fifoOut[27][11][w-1];
              unloadMuxOut[10] = fifoOut[28][11][w-1];
              unloadMuxOut[11] = fifoOut[29][11][w-1];
              unloadMuxOut[12] = fifoOut[30][11][w-1];
              unloadMuxOut[13] = fifoOut[31][11][w-1];
              unloadMuxOut[14] = fifoOut[32][11][w-1];
              unloadMuxOut[15] = fifoOut[33][11][w-1];
              unloadMuxOut[16] = fifoOut[34][11][w-1];
              unloadMuxOut[17] = fifoOut[35][11][w-1];
              unloadMuxOut[18] = fifoOut[36][11][w-1];
              unloadMuxOut[19] = fifoOut[37][11][w-1];
              unloadMuxOut[20] = fifoOut[38][11][w-1];
              unloadMuxOut[21] = fifoOut[39][11][w-1];
              unloadMuxOut[22] = fifoOut[40][11][w-1];
              unloadMuxOut[23] = fifoOut[41][11][w-1];
              unloadMuxOut[24] = fifoOut[42][11][w-1];
              unloadMuxOut[25] = fifoOut[43][11][w-1];
              unloadMuxOut[26] = fifoOut[44][11][w-1];
              unloadMuxOut[27] = fifoOut[45][11][w-1];
              unloadMuxOut[28] = fifoOut[46][11][w-1];
              unloadMuxOut[29] = fifoOut[47][11][w-1];
              unloadMuxOut[30] = fifoOut[48][11][w-1];
              unloadMuxOut[31] = fifoOut[49][11][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[50][11][w-1];
              unloadMuxOut[1] = fifoOut[51][11][w-1];
              unloadMuxOut[2] = fifoOut[26][10][w-1];
              unloadMuxOut[3] = fifoOut[27][10][w-1];
              unloadMuxOut[4] = fifoOut[28][10][w-1];
              unloadMuxOut[5] = fifoOut[29][10][w-1];
              unloadMuxOut[6] = fifoOut[30][10][w-1];
              unloadMuxOut[7] = fifoOut[31][10][w-1];
              unloadMuxOut[8] = fifoOut[32][10][w-1];
              unloadMuxOut[9] = fifoOut[33][10][w-1];
              unloadMuxOut[10] = fifoOut[34][10][w-1];
              unloadMuxOut[11] = fifoOut[35][10][w-1];
              unloadMuxOut[12] = fifoOut[36][10][w-1];
              unloadMuxOut[13] = fifoOut[37][10][w-1];
              unloadMuxOut[14] = fifoOut[38][10][w-1];
              unloadMuxOut[15] = fifoOut[39][10][w-1];
              unloadMuxOut[16] = fifoOut[40][10][w-1];
              unloadMuxOut[17] = fifoOut[41][10][w-1];
              unloadMuxOut[18] = fifoOut[42][10][w-1];
              unloadMuxOut[19] = fifoOut[43][10][w-1];
              unloadMuxOut[20] = fifoOut[44][10][w-1];
              unloadMuxOut[21] = fifoOut[45][10][w-1];
              unloadMuxOut[22] = fifoOut[46][10][w-1];
              unloadMuxOut[23] = fifoOut[47][10][w-1];
              unloadMuxOut[24] = fifoOut[48][10][w-1];
              unloadMuxOut[25] = fifoOut[49][10][w-1];
              unloadMuxOut[26] = fifoOut[50][10][w-1];
              unloadMuxOut[27] = fifoOut[51][10][w-1];
              unloadMuxOut[28] = fifoOut[26][9][w-1];
              unloadMuxOut[29] = fifoOut[27][9][w-1];
              unloadMuxOut[30] = fifoOut[28][9][w-1];
              unloadMuxOut[31] = fifoOut[29][9][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[30][9][w-1];
              unloadMuxOut[1] = fifoOut[31][9][w-1];
              unloadMuxOut[2] = fifoOut[32][9][w-1];
              unloadMuxOut[3] = fifoOut[33][9][w-1];
              unloadMuxOut[4] = fifoOut[34][9][w-1];
              unloadMuxOut[5] = fifoOut[35][9][w-1];
              unloadMuxOut[6] = fifoOut[36][9][w-1];
              unloadMuxOut[7] = fifoOut[37][9][w-1];
              unloadMuxOut[8] = fifoOut[38][9][w-1];
              unloadMuxOut[9] = fifoOut[39][9][w-1];
              unloadMuxOut[10] = fifoOut[40][9][w-1];
              unloadMuxOut[11] = fifoOut[41][9][w-1];
              unloadMuxOut[12] = fifoOut[42][9][w-1];
              unloadMuxOut[13] = fifoOut[43][9][w-1];
              unloadMuxOut[14] = fifoOut[44][9][w-1];
              unloadMuxOut[15] = fifoOut[45][9][w-1];
              unloadMuxOut[16] = fifoOut[46][9][w-1];
              unloadMuxOut[17] = fifoOut[47][9][w-1];
              unloadMuxOut[18] = fifoOut[48][9][w-1];
              unloadMuxOut[19] = fifoOut[49][9][w-1];
              unloadMuxOut[20] = fifoOut[50][9][w-1];
              unloadMuxOut[21] = fifoOut[51][9][w-1];
              unloadMuxOut[22] = fifoOut[26][8][w-1];
              unloadMuxOut[23] = fifoOut[27][8][w-1];
              unloadMuxOut[24] = fifoOut[28][8][w-1];
              unloadMuxOut[25] = fifoOut[29][8][w-1];
              unloadMuxOut[26] = fifoOut[30][8][w-1];
              unloadMuxOut[27] = fifoOut[31][8][w-1];
              unloadMuxOut[28] = fifoOut[32][8][w-1];
              unloadMuxOut[29] = fifoOut[33][8][w-1];
              unloadMuxOut[30] = fifoOut[34][8][w-1];
              unloadMuxOut[31] = fifoOut[35][8][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[36][8][w-1];
              unloadMuxOut[1] = fifoOut[37][8][w-1];
              unloadMuxOut[2] = fifoOut[38][8][w-1];
              unloadMuxOut[3] = fifoOut[39][8][w-1];
              unloadMuxOut[4] = fifoOut[40][8][w-1];
              unloadMuxOut[5] = fifoOut[41][8][w-1];
              unloadMuxOut[6] = fifoOut[42][8][w-1];
              unloadMuxOut[7] = fifoOut[43][8][w-1];
              unloadMuxOut[8] = fifoOut[44][8][w-1];
              unloadMuxOut[9] = fifoOut[45][8][w-1];
              unloadMuxOut[10] = fifoOut[46][8][w-1];
              unloadMuxOut[11] = fifoOut[47][8][w-1];
              unloadMuxOut[12] = fifoOut[48][8][w-1];
              unloadMuxOut[13] = fifoOut[49][8][w-1];
              unloadMuxOut[14] = fifoOut[50][8][w-1];
              unloadMuxOut[15] = fifoOut[51][8][w-1];
              unloadMuxOut[16] = fifoOut[26][7][w-1];
              unloadMuxOut[17] = fifoOut[27][7][w-1];
              unloadMuxOut[18] = fifoOut[28][7][w-1];
              unloadMuxOut[19] = fifoOut[29][7][w-1];
              unloadMuxOut[20] = fifoOut[30][7][w-1];
              unloadMuxOut[21] = fifoOut[31][7][w-1];
              unloadMuxOut[22] = fifoOut[32][7][w-1];
              unloadMuxOut[23] = fifoOut[33][7][w-1];
              unloadMuxOut[24] = fifoOut[34][7][w-1];
              unloadMuxOut[25] = fifoOut[35][7][w-1];
              unloadMuxOut[26] = fifoOut[36][7][w-1];
              unloadMuxOut[27] = fifoOut[37][7][w-1];
              unloadMuxOut[28] = fifoOut[38][7][w-1];
              unloadMuxOut[29] = fifoOut[39][7][w-1];
              unloadMuxOut[30] = fifoOut[40][7][w-1];
              unloadMuxOut[31] = fifoOut[41][7][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[42][7][w-1];
              unloadMuxOut[1] = fifoOut[43][7][w-1];
              unloadMuxOut[2] = fifoOut[44][7][w-1];
              unloadMuxOut[3] = fifoOut[45][7][w-1];
              unloadMuxOut[4] = fifoOut[46][7][w-1];
              unloadMuxOut[5] = fifoOut[47][7][w-1];
              unloadMuxOut[6] = fifoOut[48][7][w-1];
              unloadMuxOut[7] = fifoOut[49][7][w-1];
              unloadMuxOut[8] = fifoOut[50][7][w-1];
              unloadMuxOut[9] = fifoOut[51][7][w-1];
              unloadMuxOut[10] = fifoOut[26][6][w-1];
              unloadMuxOut[11] = fifoOut[27][6][w-1];
              unloadMuxOut[12] = fifoOut[28][6][w-1];
              unloadMuxOut[13] = fifoOut[29][6][w-1];
              unloadMuxOut[14] = fifoOut[30][6][w-1];
              unloadMuxOut[15] = fifoOut[31][6][w-1];
              unloadMuxOut[16] = fifoOut[32][6][w-1];
              unloadMuxOut[17] = fifoOut[33][6][w-1];
              unloadMuxOut[18] = fifoOut[34][6][w-1];
              unloadMuxOut[19] = fifoOut[35][6][w-1];
              unloadMuxOut[20] = fifoOut[36][6][w-1];
              unloadMuxOut[21] = fifoOut[37][6][w-1];
              unloadMuxOut[22] = fifoOut[38][6][w-1];
              unloadMuxOut[23] = fifoOut[39][6][w-1];
              unloadMuxOut[24] = fifoOut[40][6][w-1];
              unloadMuxOut[25] = fifoOut[41][6][w-1];
              unloadMuxOut[26] = fifoOut[42][6][w-1];
              unloadMuxOut[27] = fifoOut[43][6][w-1];
              unloadMuxOut[28] = fifoOut[44][6][w-1];
              unloadMuxOut[29] = fifoOut[45][6][w-1];
              unloadMuxOut[30] = fifoOut[46][6][w-1];
              unloadMuxOut[31] = fifoOut[47][6][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[48][6][w-1];
              unloadMuxOut[1] = fifoOut[49][6][w-1];
              unloadMuxOut[2] = fifoOut[50][6][w-1];
              unloadMuxOut[3] = fifoOut[51][6][w-1];
              unloadMuxOut[4] = fifoOut[26][5][w-1];
              unloadMuxOut[5] = fifoOut[27][5][w-1];
              unloadMuxOut[6] = fifoOut[28][5][w-1];
              unloadMuxOut[7] = fifoOut[29][5][w-1];
              unloadMuxOut[8] = fifoOut[30][5][w-1];
              unloadMuxOut[9] = fifoOut[31][5][w-1];
              unloadMuxOut[10] = fifoOut[32][5][w-1];
              unloadMuxOut[11] = fifoOut[33][5][w-1];
              unloadMuxOut[12] = fifoOut[34][5][w-1];
              unloadMuxOut[13] = fifoOut[35][5][w-1];
              unloadMuxOut[14] = fifoOut[36][5][w-1];
              unloadMuxOut[15] = fifoOut[37][5][w-1];
              unloadMuxOut[16] = fifoOut[38][5][w-1];
              unloadMuxOut[17] = fifoOut[39][5][w-1];
              unloadMuxOut[18] = fifoOut[40][5][w-1];
              unloadMuxOut[19] = fifoOut[41][5][w-1];
              unloadMuxOut[20] = fifoOut[42][5][w-1];
              unloadMuxOut[21] = fifoOut[43][5][w-1];
              unloadMuxOut[22] = fifoOut[44][5][w-1];
              unloadMuxOut[23] = fifoOut[45][5][w-1];
              unloadMuxOut[24] = fifoOut[46][5][w-1];
              unloadMuxOut[25] = fifoOut[47][5][w-1];
              unloadMuxOut[26] = fifoOut[48][5][w-1];
              unloadMuxOut[27] = fifoOut[49][5][w-1];
              unloadMuxOut[28] = fifoOut[50][5][w-1];
              unloadMuxOut[29] = fifoOut[51][5][w-1];
              unloadMuxOut[30] = fifoOut[26][4][w-1];
              unloadMuxOut[31] = fifoOut[27][4][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[28][4][w-1];
              unloadMuxOut[1] = fifoOut[29][4][w-1];
              unloadMuxOut[2] = fifoOut[30][4][w-1];
              unloadMuxOut[3] = fifoOut[31][4][w-1];
              unloadMuxOut[4] = fifoOut[32][4][w-1];
              unloadMuxOut[5] = fifoOut[33][4][w-1];
              unloadMuxOut[6] = fifoOut[34][4][w-1];
              unloadMuxOut[7] = fifoOut[35][4][w-1];
              unloadMuxOut[8] = fifoOut[36][4][w-1];
              unloadMuxOut[9] = fifoOut[37][4][w-1];
              unloadMuxOut[10] = fifoOut[38][4][w-1];
              unloadMuxOut[11] = fifoOut[39][4][w-1];
              unloadMuxOut[12] = fifoOut[40][4][w-1];
              unloadMuxOut[13] = fifoOut[41][4][w-1];
              unloadMuxOut[14] = fifoOut[42][4][w-1];
              unloadMuxOut[15] = fifoOut[43][4][w-1];
              unloadMuxOut[16] = fifoOut[44][4][w-1];
              unloadMuxOut[17] = fifoOut[45][4][w-1];
              unloadMuxOut[18] = fifoOut[46][4][w-1];
              unloadMuxOut[19] = fifoOut[47][4][w-1];
              unloadMuxOut[20] = fifoOut[48][4][w-1];
              unloadMuxOut[21] = fifoOut[49][4][w-1];
              unloadMuxOut[22] = fifoOut[50][4][w-1];
              unloadMuxOut[23] = fifoOut[51][4][w-1];
              unloadMuxOut[24] = fifoOut[26][3][w-1];
              unloadMuxOut[25] = fifoOut[27][3][w-1];
              unloadMuxOut[26] = fifoOut[28][3][w-1];
              unloadMuxOut[27] = fifoOut[29][3][w-1];
              unloadMuxOut[28] = fifoOut[30][3][w-1];
              unloadMuxOut[29] = fifoOut[31][3][w-1];
              unloadMuxOut[30] = fifoOut[32][3][w-1];
              unloadMuxOut[31] = fifoOut[33][3][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[34][3][w-1];
              unloadMuxOut[1] = fifoOut[35][3][w-1];
              unloadMuxOut[2] = fifoOut[36][3][w-1];
              unloadMuxOut[3] = fifoOut[37][3][w-1];
              unloadMuxOut[4] = fifoOut[38][3][w-1];
              unloadMuxOut[5] = fifoOut[39][3][w-1];
              unloadMuxOut[6] = fifoOut[40][3][w-1];
              unloadMuxOut[7] = fifoOut[41][3][w-1];
              unloadMuxOut[8] = fifoOut[42][3][w-1];
              unloadMuxOut[9] = fifoOut[43][3][w-1];
              unloadMuxOut[10] = fifoOut[44][3][w-1];
              unloadMuxOut[11] = fifoOut[45][3][w-1];
              unloadMuxOut[12] = fifoOut[46][3][w-1];
              unloadMuxOut[13] = fifoOut[47][3][w-1];
              unloadMuxOut[14] = fifoOut[48][3][w-1];
              unloadMuxOut[15] = fifoOut[49][3][w-1];
              unloadMuxOut[16] = fifoOut[50][3][w-1];
              unloadMuxOut[17] = fifoOut[51][3][w-1];
              unloadMuxOut[18] = fifoOut[26][2][w-1];
              unloadMuxOut[19] = fifoOut[27][2][w-1];
              unloadMuxOut[20] = fifoOut[28][2][w-1];
              unloadMuxOut[21] = fifoOut[29][2][w-1];
              unloadMuxOut[22] = fifoOut[30][2][w-1];
              unloadMuxOut[23] = fifoOut[31][2][w-1];
              unloadMuxOut[24] = fifoOut[32][2][w-1];
              unloadMuxOut[25] = fifoOut[33][2][w-1];
              unloadMuxOut[26] = fifoOut[34][2][w-1];
              unloadMuxOut[27] = fifoOut[35][2][w-1];
              unloadMuxOut[28] = fifoOut[36][2][w-1];
              unloadMuxOut[29] = fifoOut[37][2][w-1];
              unloadMuxOut[30] = fifoOut[38][2][w-1];
              unloadMuxOut[31] = fifoOut[39][2][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[40][2][w-1];
              unloadMuxOut[1] = fifoOut[41][2][w-1];
              unloadMuxOut[2] = fifoOut[42][2][w-1];
              unloadMuxOut[3] = fifoOut[43][2][w-1];
              unloadMuxOut[4] = fifoOut[44][2][w-1];
              unloadMuxOut[5] = fifoOut[45][2][w-1];
              unloadMuxOut[6] = fifoOut[46][2][w-1];
              unloadMuxOut[7] = fifoOut[47][2][w-1];
              unloadMuxOut[8] = fifoOut[48][2][w-1];
              unloadMuxOut[9] = fifoOut[49][2][w-1];
              unloadMuxOut[10] = fifoOut[50][2][w-1];
              unloadMuxOut[11] = fifoOut[51][2][w-1];
              unloadMuxOut[12] = fifoOut[26][1][w-1];
              unloadMuxOut[13] = fifoOut[27][1][w-1];
              unloadMuxOut[14] = fifoOut[28][1][w-1];
              unloadMuxOut[15] = fifoOut[29][1][w-1];
              unloadMuxOut[16] = fifoOut[30][1][w-1];
              unloadMuxOut[17] = fifoOut[31][1][w-1];
              unloadMuxOut[18] = fifoOut[32][1][w-1];
              unloadMuxOut[19] = fifoOut[33][1][w-1];
              unloadMuxOut[20] = fifoOut[34][1][w-1];
              unloadMuxOut[21] = fifoOut[35][1][w-1];
              unloadMuxOut[22] = fifoOut[36][1][w-1];
              unloadMuxOut[23] = fifoOut[37][1][w-1];
              unloadMuxOut[24] = fifoOut[38][1][w-1];
              unloadMuxOut[25] = fifoOut[39][1][w-1];
              unloadMuxOut[26] = fifoOut[40][1][w-1];
              unloadMuxOut[27] = fifoOut[41][1][w-1];
              unloadMuxOut[28] = fifoOut[42][1][w-1];
              unloadMuxOut[29] = fifoOut[43][1][w-1];
              unloadMuxOut[30] = fifoOut[44][1][w-1];
              unloadMuxOut[31] = fifoOut[45][1][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[46][1][w-1];
              unloadMuxOut[1] = fifoOut[47][1][w-1];
              unloadMuxOut[2] = fifoOut[48][1][w-1];
              unloadMuxOut[3] = fifoOut[49][1][w-1];
              unloadMuxOut[4] = fifoOut[50][1][w-1];
              unloadMuxOut[5] = fifoOut[51][1][w-1];
              unloadMuxOut[6] = fifoOut[26][0][w-1];
              unloadMuxOut[7] = fifoOut[27][0][w-1];
              unloadMuxOut[8] = fifoOut[28][0][w-1];
              unloadMuxOut[9] = fifoOut[29][0][w-1];
              unloadMuxOut[10] = fifoOut[0][12][w-1];
              unloadMuxOut[11] = fifoOut[1][12][w-1];
              unloadMuxOut[12] = fifoOut[2][12][w-1];
              unloadMuxOut[13] = fifoOut[3][12][w-1];
              unloadMuxOut[14] = fifoOut[4][12][w-1];
              unloadMuxOut[15] = fifoOut[5][12][w-1];
              unloadMuxOut[16] = fifoOut[6][12][w-1];
              unloadMuxOut[17] = fifoOut[7][12][w-1];
              unloadMuxOut[18] = fifoOut[8][12][w-1];
              unloadMuxOut[19] = fifoOut[9][12][w-1];
              unloadMuxOut[20] = fifoOut[10][12][w-1];
              unloadMuxOut[21] = fifoOut[11][12][w-1];
              unloadMuxOut[22] = fifoOut[12][12][w-1];
              unloadMuxOut[23] = fifoOut[13][12][w-1];
              unloadMuxOut[24] = fifoOut[14][12][w-1];
              unloadMuxOut[25] = fifoOut[15][12][w-1];
              unloadMuxOut[26] = fifoOut[16][12][w-1];
              unloadMuxOut[27] = fifoOut[17][12][w-1];
              unloadMuxOut[28] = fifoOut[18][12][w-1];
              unloadMuxOut[29] = fifoOut[19][12][w-1];
              unloadMuxOut[30] = fifoOut[20][12][w-1];
              unloadMuxOut[31] = fifoOut[21][12][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[22][12][w-1];
              unloadMuxOut[1] = fifoOut[23][12][w-1];
              unloadMuxOut[2] = fifoOut[24][12][w-1];
              unloadMuxOut[3] = fifoOut[25][12][w-1];
              unloadMuxOut[4] = fifoOut[0][11][w-1];
              unloadMuxOut[5] = fifoOut[1][11][w-1];
              unloadMuxOut[6] = fifoOut[2][11][w-1];
              unloadMuxOut[7] = fifoOut[3][11][w-1];
              unloadMuxOut[8] = fifoOut[4][11][w-1];
              unloadMuxOut[9] = fifoOut[5][11][w-1];
              unloadMuxOut[10] = fifoOut[6][11][w-1];
              unloadMuxOut[11] = fifoOut[7][11][w-1];
              unloadMuxOut[12] = fifoOut[8][11][w-1];
              unloadMuxOut[13] = fifoOut[9][11][w-1];
              unloadMuxOut[14] = fifoOut[10][11][w-1];
              unloadMuxOut[15] = fifoOut[11][11][w-1];
              unloadMuxOut[16] = fifoOut[12][11][w-1];
              unloadMuxOut[17] = fifoOut[13][11][w-1];
              unloadMuxOut[18] = fifoOut[14][11][w-1];
              unloadMuxOut[19] = fifoOut[15][11][w-1];
              unloadMuxOut[20] = fifoOut[16][11][w-1];
              unloadMuxOut[21] = fifoOut[17][11][w-1];
              unloadMuxOut[22] = fifoOut[18][11][w-1];
              unloadMuxOut[23] = fifoOut[19][11][w-1];
              unloadMuxOut[24] = fifoOut[20][11][w-1];
              unloadMuxOut[25] = fifoOut[21][11][w-1];
              unloadMuxOut[26] = fifoOut[22][11][w-1];
              unloadMuxOut[27] = fifoOut[23][11][w-1];
              unloadMuxOut[28] = fifoOut[24][11][w-1];
              unloadMuxOut[29] = fifoOut[25][11][w-1];
              unloadMuxOut[30] = fifoOut[0][10][w-1];
              unloadMuxOut[31] = fifoOut[1][10][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[2][10][w-1];
              unloadMuxOut[1] = fifoOut[3][10][w-1];
              unloadMuxOut[2] = fifoOut[4][10][w-1];
              unloadMuxOut[3] = fifoOut[5][10][w-1];
              unloadMuxOut[4] = fifoOut[6][10][w-1];
              unloadMuxOut[5] = fifoOut[7][10][w-1];
              unloadMuxOut[6] = fifoOut[8][10][w-1];
              unloadMuxOut[7] = fifoOut[9][10][w-1];
              unloadMuxOut[8] = fifoOut[10][10][w-1];
              unloadMuxOut[9] = fifoOut[11][10][w-1];
              unloadMuxOut[10] = fifoOut[12][10][w-1];
              unloadMuxOut[11] = fifoOut[13][10][w-1];
              unloadMuxOut[12] = fifoOut[14][10][w-1];
              unloadMuxOut[13] = fifoOut[15][10][w-1];
              unloadMuxOut[14] = fifoOut[16][10][w-1];
              unloadMuxOut[15] = fifoOut[17][10][w-1];
              unloadMuxOut[16] = fifoOut[18][10][w-1];
              unloadMuxOut[17] = fifoOut[19][10][w-1];
              unloadMuxOut[18] = fifoOut[20][10][w-1];
              unloadMuxOut[19] = fifoOut[21][10][w-1];
              unloadMuxOut[20] = fifoOut[22][10][w-1];
              unloadMuxOut[21] = fifoOut[23][10][w-1];
              unloadMuxOut[22] = fifoOut[24][10][w-1];
              unloadMuxOut[23] = fifoOut[25][10][w-1];
              unloadMuxOut[24] = fifoOut[0][9][w-1];
              unloadMuxOut[25] = fifoOut[1][9][w-1];
              unloadMuxOut[26] = fifoOut[2][9][w-1];
              unloadMuxOut[27] = fifoOut[3][9][w-1];
              unloadMuxOut[28] = fifoOut[4][9][w-1];
              unloadMuxOut[29] = fifoOut[5][9][w-1];
              unloadMuxOut[30] = fifoOut[6][9][w-1];
              unloadMuxOut[31] = fifoOut[7][9][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[8][9][w-1];
              unloadMuxOut[1] = fifoOut[9][9][w-1];
              unloadMuxOut[2] = fifoOut[10][9][w-1];
              unloadMuxOut[3] = fifoOut[11][9][w-1];
              unloadMuxOut[4] = fifoOut[12][9][w-1];
              unloadMuxOut[5] = fifoOut[13][9][w-1];
              unloadMuxOut[6] = fifoOut[14][9][w-1];
              unloadMuxOut[7] = fifoOut[15][9][w-1];
              unloadMuxOut[8] = fifoOut[16][9][w-1];
              unloadMuxOut[9] = fifoOut[17][9][w-1];
              unloadMuxOut[10] = fifoOut[18][9][w-1];
              unloadMuxOut[11] = fifoOut[19][9][w-1];
              unloadMuxOut[12] = fifoOut[20][9][w-1];
              unloadMuxOut[13] = fifoOut[21][9][w-1];
              unloadMuxOut[14] = fifoOut[22][9][w-1];
              unloadMuxOut[15] = fifoOut[23][9][w-1];
              unloadMuxOut[16] = fifoOut[24][9][w-1];
              unloadMuxOut[17] = fifoOut[25][9][w-1];
              unloadMuxOut[18] = fifoOut[0][8][w-1];
              unloadMuxOut[19] = fifoOut[1][8][w-1];
              unloadMuxOut[20] = fifoOut[2][8][w-1];
              unloadMuxOut[21] = fifoOut[3][8][w-1];
              unloadMuxOut[22] = fifoOut[4][8][w-1];
              unloadMuxOut[23] = fifoOut[5][8][w-1];
              unloadMuxOut[24] = fifoOut[6][8][w-1];
              unloadMuxOut[25] = fifoOut[7][8][w-1];
              unloadMuxOut[26] = fifoOut[8][8][w-1];
              unloadMuxOut[27] = fifoOut[9][8][w-1];
              unloadMuxOut[28] = fifoOut[10][8][w-1];
              unloadMuxOut[29] = fifoOut[11][8][w-1];
              unloadMuxOut[30] = fifoOut[12][8][w-1];
              unloadMuxOut[31] = fifoOut[13][8][w-1];
       end
       16: begin
              unloadMuxOut[0] = fifoOut[14][8][w-1];
              unloadMuxOut[1] = fifoOut[15][8][w-1];
              unloadMuxOut[2] = fifoOut[16][8][w-1];
              unloadMuxOut[3] = fifoOut[17][8][w-1];
              unloadMuxOut[4] = fifoOut[18][8][w-1];
              unloadMuxOut[5] = fifoOut[19][8][w-1];
              unloadMuxOut[6] = fifoOut[20][8][w-1];
              unloadMuxOut[7] = fifoOut[21][8][w-1];
              unloadMuxOut[8] = fifoOut[22][8][w-1];
              unloadMuxOut[9] = fifoOut[23][8][w-1];
              unloadMuxOut[10] = fifoOut[24][8][w-1];
              unloadMuxOut[11] = fifoOut[25][8][w-1];
              unloadMuxOut[12] = fifoOut[0][7][w-1];
              unloadMuxOut[13] = fifoOut[1][7][w-1];
              unloadMuxOut[14] = fifoOut[2][7][w-1];
              unloadMuxOut[15] = fifoOut[3][7][w-1];
              unloadMuxOut[16] = fifoOut[4][7][w-1];
              unloadMuxOut[17] = fifoOut[5][7][w-1];
              unloadMuxOut[18] = fifoOut[6][7][w-1];
              unloadMuxOut[19] = fifoOut[7][7][w-1];
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0;
             end
       end
    endcase
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[0][6];
              muxOutConnector[1] = fifoOut[1][6];
              muxOutConnector[2] = fifoOut[2][6];
              muxOutConnector[3] = fifoOut[3][6];
              muxOutConnector[4] = fifoOut[4][6];
              muxOutConnector[5] = fifoOut[5][6];
              muxOutConnector[6] = fifoOut[6][6];
              muxOutConnector[7] = fifoOut[7][6];
              muxOutConnector[8] = fifoOut[8][6];
              muxOutConnector[9] = fifoOut[9][6];
              muxOutConnector[10] = fifoOut[10][6];
              muxOutConnector[11] = fifoOut[11][6];
              muxOutConnector[12] = fifoOut[12][6];
              muxOutConnector[13] = fifoOut[13][6];
              muxOutConnector[14] = fifoOut[14][6];
              muxOutConnector[15] = fifoOut[15][6];
              muxOutConnector[16] = fifoOut[16][6];
              muxOutConnector[17] = fifoOut[17][6];
              muxOutConnector[18] = fifoOut[18][6];
              muxOutConnector[19] = fifoOut[19][6];
              muxOutConnector[20] = fifoOut[20][6];
              muxOutConnector[21] = fifoOut[21][6];
              muxOutConnector[22] = fifoOut[22][6];
              muxOutConnector[23] = fifoOut[23][6];
              muxOutConnector[24] = fifoOut[24][6];
              muxOutConnector[25] = fifoOut[25][6];
              muxOutConnector[26] = fifoOut[42][4];
              muxOutConnector[27] = fifoOut[43][4];
              muxOutConnector[28] = fifoOut[44][4];
              muxOutConnector[29] = fifoOut[45][4];
              muxOutConnector[30] = fifoOut[46][4];
              muxOutConnector[31] = fifoOut[47][4];
              muxOutConnector[32] = fifoOut[48][4];
              muxOutConnector[33] = fifoOut[49][4];
              muxOutConnector[34] = fifoOut[50][4];
              muxOutConnector[35] = fifoOut[51][4];
              muxOutConnector[36] = fifoOut[26][3];
              muxOutConnector[37] = fifoOut[27][3];
              muxOutConnector[38] = fifoOut[28][3];
              muxOutConnector[39] = fifoOut[29][3];
              muxOutConnector[40] = fifoOut[30][3];
              muxOutConnector[41] = fifoOut[31][3];
              muxOutConnector[42] = fifoOut[32][3];
              muxOutConnector[43] = fifoOut[33][3];
              muxOutConnector[44] = fifoOut[34][3];
              muxOutConnector[45] = fifoOut[35][3];
              muxOutConnector[46] = fifoOut[36][3];
              muxOutConnector[47] = fifoOut[37][3];
              muxOutConnector[48] = fifoOut[38][3];
              muxOutConnector[49] = fifoOut[39][3];
              muxOutConnector[50] = fifoOut[40][3];
              muxOutConnector[51] = fifoOut[41][3];
       end
       1: begin
              muxOutConnector[0] = fifoOut[0][6];
              muxOutConnector[1] = fifoOut[1][6];
              muxOutConnector[2] = fifoOut[2][6];
              muxOutConnector[3] = fifoOut[3][6];
              muxOutConnector[4] = fifoOut[4][6];
              muxOutConnector[5] = fifoOut[5][6];
              muxOutConnector[6] = fifoOut[6][6];
              muxOutConnector[7] = fifoOut[7][6];
              muxOutConnector[8] = fifoOut[8][6];
              muxOutConnector[9] = fifoOut[9][6];
              muxOutConnector[10] = fifoOut[10][6];
              muxOutConnector[11] = fifoOut[11][6];
              muxOutConnector[12] = fifoOut[12][6];
              muxOutConnector[13] = fifoOut[13][6];
              muxOutConnector[14] = fifoOut[14][6];
              muxOutConnector[15] = fifoOut[15][6];
              muxOutConnector[16] = fifoOut[16][6];
              muxOutConnector[17] = fifoOut[17][6];
              muxOutConnector[18] = fifoOut[18][6];
              muxOutConnector[19] = fifoOut[19][6];
              muxOutConnector[20] = fifoOut[20][6];
              muxOutConnector[21] = fifoOut[21][6];
              muxOutConnector[22] = fifoOut[22][6];
              muxOutConnector[23] = fifoOut[23][6];
              muxOutConnector[24] = fifoOut[24][6];
              muxOutConnector[25] = fifoOut[25][6];
              muxOutConnector[26] = fifoOut[42][4];
              muxOutConnector[27] = fifoOut[43][4];
              muxOutConnector[28] = fifoOut[44][4];
              muxOutConnector[29] = fifoOut[45][4];
              muxOutConnector[30] = fifoOut[46][4];
              muxOutConnector[31] = fifoOut[47][4];
              muxOutConnector[32] = fifoOut[48][4];
              muxOutConnector[33] = fifoOut[49][4];
              muxOutConnector[34] = fifoOut[50][4];
              muxOutConnector[35] = fifoOut[51][4];
              muxOutConnector[36] = fifoOut[26][3];
              muxOutConnector[37] = fifoOut[27][3];
              muxOutConnector[38] = fifoOut[28][3];
              muxOutConnector[39] = fifoOut[29][3];
              muxOutConnector[40] = fifoOut[30][3];
              muxOutConnector[41] = fifoOut[31][3];
              muxOutConnector[42] = fifoOut[32][3];
              muxOutConnector[43] = fifoOut[33][3];
              muxOutConnector[44] = fifoOut[34][3];
              muxOutConnector[45] = fifoOut[35][3];
              muxOutConnector[46] = fifoOut[36][3];
              muxOutConnector[47] = fifoOut[37][3];
              muxOutConnector[48] = fifoOut[38][3];
              muxOutConnector[49] = fifoOut[39][3];
              muxOutConnector[50] = fifoOut[40][3];
              muxOutConnector[51] = fifoOut[41][3];
       end
       2: begin
              muxOutConnector[0] = fifoOut[0][6];
              muxOutConnector[1] = fifoOut[1][6];
              muxOutConnector[2] = fifoOut[2][6];
              muxOutConnector[3] = fifoOut[3][6];
              muxOutConnector[4] = fifoOut[4][6];
              muxOutConnector[5] = fifoOut[5][6];
              muxOutConnector[6] = fifoOut[6][6];
              muxOutConnector[7] = fifoOut[7][6];
              muxOutConnector[8] = fifoOut[8][6];
              muxOutConnector[9] = fifoOut[9][6];
              muxOutConnector[10] = fifoOut[10][6];
              muxOutConnector[11] = fifoOut[11][6];
              muxOutConnector[12] = fifoOut[12][6];
              muxOutConnector[13] = fifoOut[13][6];
              muxOutConnector[14] = fifoOut[14][6];
              muxOutConnector[15] = fifoOut[15][6];
              muxOutConnector[16] = fifoOut[16][6];
              muxOutConnector[17] = fifoOut[17][6];
              muxOutConnector[18] = fifoOut[18][6];
              muxOutConnector[19] = fifoOut[19][6];
              muxOutConnector[20] = fifoOut[20][6];
              muxOutConnector[21] = fifoOut[21][6];
              muxOutConnector[22] = fifoOut[22][6];
              muxOutConnector[23] = fifoOut[23][6];
              muxOutConnector[24] = fifoOut[24][6];
              muxOutConnector[25] = fifoOut[25][6];
              muxOutConnector[26] = fifoOut[42][4];
              muxOutConnector[27] = fifoOut[43][4];
              muxOutConnector[28] = fifoOut[44][4];
              muxOutConnector[29] = fifoOut[45][4];
              muxOutConnector[30] = fifoOut[46][4];
              muxOutConnector[31] = fifoOut[47][4];
              muxOutConnector[32] = fifoOut[48][4];
              muxOutConnector[33] = fifoOut[49][4];
              muxOutConnector[34] = fifoOut[50][4];
              muxOutConnector[35] = fifoOut[51][4];
              muxOutConnector[36] = fifoOut[26][3];
              muxOutConnector[37] = fifoOut[27][3];
              muxOutConnector[38] = fifoOut[28][3];
              muxOutConnector[39] = fifoOut[29][3];
              muxOutConnector[40] = fifoOut[30][3];
              muxOutConnector[41] = fifoOut[31][3];
              muxOutConnector[42] = fifoOut[32][3];
              muxOutConnector[43] = fifoOut[33][3];
              muxOutConnector[44] = fifoOut[34][3];
              muxOutConnector[45] = fifoOut[35][3];
              muxOutConnector[46] = fifoOut[36][3];
              muxOutConnector[47] = fifoOut[37][3];
              muxOutConnector[48] = fifoOut[38][3];
              muxOutConnector[49] = fifoOut[39][3];
              muxOutConnector[50] = fifoOut[40][3];
              muxOutConnector[51] = fifoOut[41][3];
       end
       3: begin
              muxOutConnector[0] = fifoOut[0][6];
              muxOutConnector[1] = fifoOut[1][6];
              muxOutConnector[2] = fifoOut[2][6];
              muxOutConnector[3] = fifoOut[3][6];
              muxOutConnector[4] = fifoOut[4][6];
              muxOutConnector[5] = fifoOut[5][6];
              muxOutConnector[6] = fifoOut[6][6];
              muxOutConnector[7] = fifoOut[7][6];
              muxOutConnector[8] = fifoOut[8][6];
              muxOutConnector[9] = fifoOut[9][6];
              muxOutConnector[10] = fifoOut[10][6];
              muxOutConnector[11] = fifoOut[11][6];
              muxOutConnector[12] = fifoOut[12][6];
              muxOutConnector[13] = fifoOut[13][6];
              muxOutConnector[14] = fifoOut[14][6];
              muxOutConnector[15] = fifoOut[15][6];
              muxOutConnector[16] = fifoOut[16][6];
              muxOutConnector[17] = fifoOut[17][6];
              muxOutConnector[18] = fifoOut[18][6];
              muxOutConnector[19] = fifoOut[19][6];
              muxOutConnector[20] = fifoOut[20][6];
              muxOutConnector[21] = fifoOut[21][6];
              muxOutConnector[22] = fifoOut[22][6];
              muxOutConnector[23] = fifoOut[23][6];
              muxOutConnector[24] = fifoOut[24][6];
              muxOutConnector[25] = fifoOut[25][6];
              muxOutConnector[26] = fifoOut[42][4];
              muxOutConnector[27] = fifoOut[43][4];
              muxOutConnector[28] = fifoOut[44][4];
              muxOutConnector[29] = fifoOut[45][4];
              muxOutConnector[30] = fifoOut[46][4];
              muxOutConnector[31] = fifoOut[47][4];
              muxOutConnector[32] = fifoOut[48][4];
              muxOutConnector[33] = fifoOut[49][4];
              muxOutConnector[34] = fifoOut[50][4];
              muxOutConnector[35] = fifoOut[51][4];
              muxOutConnector[36] = fifoOut[26][3];
              muxOutConnector[37] = fifoOut[27][3];
              muxOutConnector[38] = fifoOut[28][3];
              muxOutConnector[39] = fifoOut[29][3];
              muxOutConnector[40] = fifoOut[30][3];
              muxOutConnector[41] = fifoOut[31][3];
              muxOutConnector[42] = fifoOut[32][3];
              muxOutConnector[43] = fifoOut[33][3];
              muxOutConnector[44] = fifoOut[34][3];
              muxOutConnector[45] = fifoOut[35][3];
              muxOutConnector[46] = fifoOut[36][3];
              muxOutConnector[47] = fifoOut[37][3];
              muxOutConnector[48] = fifoOut[38][3];
              muxOutConnector[49] = fifoOut[39][3];
              muxOutConnector[50] = fifoOut[40][3];
              muxOutConnector[51] = fifoOut[41][3];
       end
       4: begin
              muxOutConnector[0] = fifoOut[0][6];
              muxOutConnector[1] = fifoOut[1][6];
              muxOutConnector[2] = fifoOut[2][6];
              muxOutConnector[3] = fifoOut[3][6];
              muxOutConnector[4] = fifoOut[4][6];
              muxOutConnector[5] = fifoOut[5][6];
              muxOutConnector[6] = fifoOut[6][6];
              muxOutConnector[7] = fifoOut[7][6];
              muxOutConnector[8] = fifoOut[8][6];
              muxOutConnector[9] = fifoOut[9][6];
              muxOutConnector[10] = fifoOut[10][6];
              muxOutConnector[11] = fifoOut[11][6];
              muxOutConnector[12] = fifoOut[12][6];
              muxOutConnector[13] = fifoOut[13][6];
              muxOutConnector[14] = fifoOut[14][6];
              muxOutConnector[15] = fifoOut[15][6];
              muxOutConnector[16] = fifoOut[16][6];
              muxOutConnector[17] = fifoOut[17][6];
              muxOutConnector[18] = fifoOut[18][6];
              muxOutConnector[19] = fifoOut[19][6];
              muxOutConnector[20] = fifoOut[20][6];
              muxOutConnector[21] = fifoOut[21][6];
              muxOutConnector[22] = fifoOut[22][6];
              muxOutConnector[23] = fifoOut[23][6];
              muxOutConnector[24] = fifoOut[24][6];
              muxOutConnector[25] = fifoOut[25][6];
              muxOutConnector[26] = fifoOut[42][4];
              muxOutConnector[27] = fifoOut[13][3];
              muxOutConnector[28] = fifoOut[14][3];
              muxOutConnector[29] = fifoOut[15][3];
              muxOutConnector[30] = fifoOut[16][3];
              muxOutConnector[31] = fifoOut[17][3];
              muxOutConnector[32] = fifoOut[18][3];
              muxOutConnector[33] = fifoOut[19][3];
              muxOutConnector[34] = fifoOut[20][3];
              muxOutConnector[35] = fifoOut[21][3];
              muxOutConnector[36] = fifoOut[22][3];
              muxOutConnector[37] = fifoOut[23][3];
              muxOutConnector[38] = fifoOut[24][3];
              muxOutConnector[39] = fifoOut[25][3];
              muxOutConnector[40] = fifoOut[0][2];
              muxOutConnector[41] = fifoOut[1][2];
              muxOutConnector[42] = fifoOut[2][2];
              muxOutConnector[43] = fifoOut[3][2];
              muxOutConnector[44] = fifoOut[4][2];
              muxOutConnector[45] = fifoOut[5][2];
              muxOutConnector[46] = fifoOut[6][2];
              muxOutConnector[47] = fifoOut[7][2];
              muxOutConnector[48] = fifoOut[8][2];
              muxOutConnector[49] = fifoOut[9][2];
              muxOutConnector[50] = fifoOut[10][2];
              muxOutConnector[51] = fifoOut[11][2];
       end
       5: begin
              muxOutConnector[0] = fifoOut[0][6];
              muxOutConnector[1] = fifoOut[1][6];
              muxOutConnector[2] = fifoOut[2][6];
              muxOutConnector[3] = fifoOut[3][6];
              muxOutConnector[4] = fifoOut[4][6];
              muxOutConnector[5] = fifoOut[5][6];
              muxOutConnector[6] = fifoOut[6][6];
              muxOutConnector[7] = fifoOut[7][6];
              muxOutConnector[8] = fifoOut[8][6];
              muxOutConnector[9] = fifoOut[9][6];
              muxOutConnector[10] = fifoOut[10][6];
              muxOutConnector[11] = fifoOut[11][6];
              muxOutConnector[12] = fifoOut[12][6];
              muxOutConnector[13] = fifoOut[13][6];
              muxOutConnector[14] = fifoOut[14][6];
              muxOutConnector[15] = fifoOut[15][6];
              muxOutConnector[16] = fifoOut[16][6];
              muxOutConnector[17] = fifoOut[17][6];
              muxOutConnector[18] = fifoOut[18][6];
              muxOutConnector[19] = fifoOut[19][6];
              muxOutConnector[20] = fifoOut[20][6];
              muxOutConnector[21] = fifoOut[21][6];
              muxOutConnector[22] = fifoOut[22][6];
              muxOutConnector[23] = fifoOut[23][6];
              muxOutConnector[24] = fifoOut[24][6];
              muxOutConnector[25] = fifoOut[25][6];
              muxOutConnector[26] = fifoOut[12][3];
              muxOutConnector[27] = fifoOut[13][3];
              muxOutConnector[28] = fifoOut[14][3];
              muxOutConnector[29] = fifoOut[15][3];
              muxOutConnector[30] = fifoOut[16][3];
              muxOutConnector[31] = fifoOut[17][3];
              muxOutConnector[32] = fifoOut[18][3];
              muxOutConnector[33] = fifoOut[19][3];
              muxOutConnector[34] = fifoOut[20][3];
              muxOutConnector[35] = fifoOut[21][3];
              muxOutConnector[36] = fifoOut[22][3];
              muxOutConnector[37] = fifoOut[23][3];
              muxOutConnector[38] = fifoOut[24][3];
              muxOutConnector[39] = fifoOut[25][3];
              muxOutConnector[40] = fifoOut[0][2];
              muxOutConnector[41] = fifoOut[1][2];
              muxOutConnector[42] = fifoOut[2][2];
              muxOutConnector[43] = fifoOut[3][2];
              muxOutConnector[44] = fifoOut[4][2];
              muxOutConnector[45] = fifoOut[5][2];
              muxOutConnector[46] = fifoOut[6][2];
              muxOutConnector[47] = fifoOut[7][2];
              muxOutConnector[48] = fifoOut[8][2];
              muxOutConnector[49] = fifoOut[9][2];
              muxOutConnector[50] = fifoOut[10][2];
              muxOutConnector[51] = fifoOut[11][2];
       end
       6: begin
              muxOutConnector[0] = fifoOut[0][6];
              muxOutConnector[1] = fifoOut[1][6];
              muxOutConnector[2] = fifoOut[2][6];
              muxOutConnector[3] = fifoOut[3][6];
              muxOutConnector[4] = fifoOut[4][6];
              muxOutConnector[5] = fifoOut[5][6];
              muxOutConnector[6] = fifoOut[6][6];
              muxOutConnector[7] = fifoOut[7][6];
              muxOutConnector[8] = fifoOut[8][6];
              muxOutConnector[9] = fifoOut[9][6];
              muxOutConnector[10] = fifoOut[10][6];
              muxOutConnector[11] = fifoOut[11][6];
              muxOutConnector[12] = fifoOut[12][6];
              muxOutConnector[13] = fifoOut[13][6];
              muxOutConnector[14] = fifoOut[14][6];
              muxOutConnector[15] = fifoOut[15][6];
              muxOutConnector[16] = fifoOut[16][6];
              muxOutConnector[17] = fifoOut[30][0];
              muxOutConnector[18] = fifoOut[31][0];
              muxOutConnector[19] = fifoOut[32][0];
              muxOutConnector[20] = fifoOut[33][0];
              muxOutConnector[21] = fifoOut[34][0];
              muxOutConnector[22] = fifoOut[35][0];
              muxOutConnector[23] = fifoOut[36][0];
              muxOutConnector[24] = fifoOut[37][0];
              muxOutConnector[25] = fifoOut[38][0];
              muxOutConnector[26] = fifoOut[12][3];
              muxOutConnector[27] = fifoOut[13][3];
              muxOutConnector[28] = fifoOut[14][3];
              muxOutConnector[29] = fifoOut[15][3];
              muxOutConnector[30] = fifoOut[16][3];
              muxOutConnector[31] = fifoOut[17][3];
              muxOutConnector[32] = fifoOut[18][3];
              muxOutConnector[33] = fifoOut[19][3];
              muxOutConnector[34] = fifoOut[20][3];
              muxOutConnector[35] = fifoOut[21][3];
              muxOutConnector[36] = fifoOut[22][3];
              muxOutConnector[37] = fifoOut[23][3];
              muxOutConnector[38] = fifoOut[24][3];
              muxOutConnector[39] = fifoOut[25][3];
              muxOutConnector[40] = fifoOut[0][2];
              muxOutConnector[41] = fifoOut[1][2];
              muxOutConnector[42] = fifoOut[2][2];
              muxOutConnector[43] = fifoOut[3][2];
              muxOutConnector[44] = fifoOut[4][2];
              muxOutConnector[45] = fifoOut[5][2];
              muxOutConnector[46] = fifoOut[6][2];
              muxOutConnector[47] = fifoOut[7][2];
              muxOutConnector[48] = fifoOut[8][2];
              muxOutConnector[49] = fifoOut[9][2];
              muxOutConnector[50] = fifoOut[10][2];
              muxOutConnector[51] = fifoOut[11][2];
       end
       7: begin
              muxOutConnector[0] = fifoOut[39][1];
              muxOutConnector[1] = fifoOut[40][1];
              muxOutConnector[2] = fifoOut[41][1];
              muxOutConnector[3] = fifoOut[42][1];
              muxOutConnector[4] = fifoOut[43][1];
              muxOutConnector[5] = fifoOut[44][1];
              muxOutConnector[6] = fifoOut[45][1];
              muxOutConnector[7] = fifoOut[46][1];
              muxOutConnector[8] = fifoOut[47][1];
              muxOutConnector[9] = fifoOut[48][1];
              muxOutConnector[10] = fifoOut[49][1];
              muxOutConnector[11] = fifoOut[50][1];
              muxOutConnector[12] = fifoOut[51][1];
              muxOutConnector[13] = fifoOut[26][0];
              muxOutConnector[14] = fifoOut[27][0];
              muxOutConnector[15] = fifoOut[28][0];
              muxOutConnector[16] = fifoOut[29][0];
              muxOutConnector[17] = fifoOut[30][0];
              muxOutConnector[18] = fifoOut[31][0];
              muxOutConnector[19] = fifoOut[32][0];
              muxOutConnector[20] = fifoOut[33][0];
              muxOutConnector[21] = fifoOut[34][0];
              muxOutConnector[22] = fifoOut[35][0];
              muxOutConnector[23] = fifoOut[36][0];
              muxOutConnector[24] = fifoOut[37][0];
              muxOutConnector[25] = fifoOut[38][0];
              muxOutConnector[26] = fifoOut[12][3];
              muxOutConnector[27] = fifoOut[13][3];
              muxOutConnector[28] = fifoOut[14][3];
              muxOutConnector[29] = fifoOut[15][3];
              muxOutConnector[30] = fifoOut[16][3];
              muxOutConnector[31] = fifoOut[17][3];
              muxOutConnector[32] = fifoOut[18][3];
              muxOutConnector[33] = fifoOut[19][3];
              muxOutConnector[34] = fifoOut[20][3];
              muxOutConnector[35] = fifoOut[21][3];
              muxOutConnector[36] = fifoOut[22][3];
              muxOutConnector[37] = fifoOut[23][3];
              muxOutConnector[38] = fifoOut[24][3];
              muxOutConnector[39] = fifoOut[25][3];
              muxOutConnector[40] = fifoOut[0][2];
              muxOutConnector[41] = fifoOut[1][2];
              muxOutConnector[42] = fifoOut[2][2];
              muxOutConnector[43] = fifoOut[3][2];
              muxOutConnector[44] = fifoOut[4][2];
              muxOutConnector[45] = fifoOut[5][2];
              muxOutConnector[46] = fifoOut[6][2];
              muxOutConnector[47] = fifoOut[7][2];
              muxOutConnector[48] = fifoOut[8][2];
              muxOutConnector[49] = fifoOut[9][2];
              muxOutConnector[50] = fifoOut[10][2];
              muxOutConnector[51] = fifoOut[11][2];
       end
       8: begin
              muxOutConnector[0] = fifoOut[39][1];
              muxOutConnector[1] = fifoOut[40][1];
              muxOutConnector[2] = fifoOut[41][1];
              muxOutConnector[3] = fifoOut[42][1];
              muxOutConnector[4] = fifoOut[43][1];
              muxOutConnector[5] = fifoOut[44][1];
              muxOutConnector[6] = fifoOut[45][1];
              muxOutConnector[7] = fifoOut[46][1];
              muxOutConnector[8] = fifoOut[47][1];
              muxOutConnector[9] = fifoOut[48][1];
              muxOutConnector[10] = fifoOut[49][1];
              muxOutConnector[11] = fifoOut[50][1];
              muxOutConnector[12] = fifoOut[51][1];
              muxOutConnector[13] = fifoOut[26][0];
              muxOutConnector[14] = fifoOut[27][0];
              muxOutConnector[15] = fifoOut[28][0];
              muxOutConnector[16] = fifoOut[29][0];
              muxOutConnector[17] = fifoOut[30][0];
              muxOutConnector[18] = fifoOut[31][0];
              muxOutConnector[19] = fifoOut[32][0];
              muxOutConnector[20] = fifoOut[33][0];
              muxOutConnector[21] = fifoOut[34][0];
              muxOutConnector[22] = fifoOut[35][0];
              muxOutConnector[23] = fifoOut[36][0];
              muxOutConnector[24] = fifoOut[37][0];
              muxOutConnector[25] = fifoOut[38][0];
              muxOutConnector[26] = fifoOut[12][3];
              muxOutConnector[27] = fifoOut[13][3];
              muxOutConnector[28] = fifoOut[14][3];
              muxOutConnector[29] = fifoOut[15][3];
              muxOutConnector[30] = fifoOut[16][3];
              muxOutConnector[31] = fifoOut[17][3];
              muxOutConnector[32] = fifoOut[18][3];
              muxOutConnector[33] = fifoOut[19][3];
              muxOutConnector[34] = fifoOut[20][3];
              muxOutConnector[35] = fifoOut[21][3];
              muxOutConnector[36] = fifoOut[22][3];
              muxOutConnector[37] = fifoOut[23][3];
              muxOutConnector[38] = fifoOut[24][3];
              muxOutConnector[39] = fifoOut[25][3];
              muxOutConnector[40] = fifoOut[0][2];
              muxOutConnector[41] = fifoOut[1][2];
              muxOutConnector[42] = fifoOut[2][2];
              muxOutConnector[43] = fifoOut[3][2];
              muxOutConnector[44] = fifoOut[4][2];
              muxOutConnector[45] = fifoOut[5][2];
              muxOutConnector[46] = fifoOut[6][2];
              muxOutConnector[47] = fifoOut[7][2];
              muxOutConnector[48] = fifoOut[8][2];
              muxOutConnector[49] = fifoOut[9][2];
              muxOutConnector[50] = fifoOut[10][2];
              muxOutConnector[51] = fifoOut[11][2];
       end
       9: begin
              muxOutConnector[0] = fifoOut[39][1];
              muxOutConnector[1] = fifoOut[40][1];
              muxOutConnector[2] = fifoOut[41][1];
              muxOutConnector[3] = fifoOut[42][1];
              muxOutConnector[4] = fifoOut[43][1];
              muxOutConnector[5] = fifoOut[44][1];
              muxOutConnector[6] = fifoOut[45][1];
              muxOutConnector[7] = fifoOut[46][1];
              muxOutConnector[8] = fifoOut[47][1];
              muxOutConnector[9] = fifoOut[48][1];
              muxOutConnector[10] = fifoOut[49][1];
              muxOutConnector[11] = fifoOut[50][1];
              muxOutConnector[12] = fifoOut[51][1];
              muxOutConnector[13] = fifoOut[26][0];
              muxOutConnector[14] = fifoOut[27][0];
              muxOutConnector[15] = fifoOut[28][0];
              muxOutConnector[16] = fifoOut[29][0];
              muxOutConnector[17] = fifoOut[30][0];
              muxOutConnector[18] = fifoOut[31][0];
              muxOutConnector[19] = fifoOut[32][0];
              muxOutConnector[20] = fifoOut[33][0];
              muxOutConnector[21] = fifoOut[34][0];
              muxOutConnector[22] = fifoOut[35][0];
              muxOutConnector[23] = fifoOut[36][0];
              muxOutConnector[24] = fifoOut[37][0];
              muxOutConnector[25] = fifoOut[38][0];
              muxOutConnector[26] = fifoOut[12][3];
              muxOutConnector[27] = fifoOut[13][3];
              muxOutConnector[28] = fifoOut[14][3];
              muxOutConnector[29] = fifoOut[15][3];
              muxOutConnector[30] = fifoOut[16][3];
              muxOutConnector[31] = fifoOut[17][3];
              muxOutConnector[32] = fifoOut[18][3];
              muxOutConnector[33] = fifoOut[19][3];
              muxOutConnector[34] = fifoOut[20][3];
              muxOutConnector[35] = fifoOut[21][3];
              muxOutConnector[36] = fifoOut[22][3];
              muxOutConnector[37] = fifoOut[23][3];
              muxOutConnector[38] = fifoOut[24][3];
              muxOutConnector[39] = fifoOut[25][3];
              muxOutConnector[40] = fifoOut[0][2];
              muxOutConnector[41] = fifoOut[1][2];
              muxOutConnector[42] = fifoOut[2][2];
              muxOutConnector[43] = fifoOut[3][2];
              muxOutConnector[44] = fifoOut[4][2];
              muxOutConnector[45] = fifoOut[5][2];
              muxOutConnector[46] = fifoOut[6][2];
              muxOutConnector[47] = fifoOut[7][2];
              muxOutConnector[48] = fifoOut[8][2];
              muxOutConnector[49] = fifoOut[9][2];
              muxOutConnector[50] = fifoOut[10][2];
              muxOutConnector[51] = fifoOut[11][2];
       end
       10: begin
              muxOutConnector[0] = fifoOut[39][1];
              muxOutConnector[1] = fifoOut[40][1];
              muxOutConnector[2] = fifoOut[41][1];
              muxOutConnector[3] = fifoOut[42][1];
              muxOutConnector[4] = fifoOut[43][1];
              muxOutConnector[5] = fifoOut[44][1];
              muxOutConnector[6] = fifoOut[45][1];
              muxOutConnector[7] = fifoOut[46][1];
              muxOutConnector[8] = fifoOut[47][1];
              muxOutConnector[9] = fifoOut[48][1];
              muxOutConnector[10] = fifoOut[49][1];
              muxOutConnector[11] = fifoOut[50][1];
              muxOutConnector[12] = fifoOut[51][1];
              muxOutConnector[13] = fifoOut[26][0];
              muxOutConnector[14] = fifoOut[27][0];
              muxOutConnector[15] = fifoOut[28][0];
              muxOutConnector[16] = fifoOut[29][0];
              muxOutConnector[17] = fifoOut[30][0];
              muxOutConnector[18] = fifoOut[31][0];
              muxOutConnector[19] = fifoOut[32][0];
              muxOutConnector[20] = fifoOut[33][0];
              muxOutConnector[21] = fifoOut[34][0];
              muxOutConnector[22] = fifoOut[35][0];
              muxOutConnector[23] = fifoOut[36][0];
              muxOutConnector[24] = fifoOut[37][0];
              muxOutConnector[25] = fifoOut[38][0];
              muxOutConnector[26] = fifoOut[12][3];
              muxOutConnector[27] = fifoOut[13][3];
              muxOutConnector[28] = fifoOut[14][3];
              muxOutConnector[29] = fifoOut[15][3];
              muxOutConnector[30] = fifoOut[16][3];
              muxOutConnector[31] = fifoOut[17][3];
              muxOutConnector[32] = fifoOut[18][3];
              muxOutConnector[33] = fifoOut[19][3];
              muxOutConnector[34] = fifoOut[20][3];
              muxOutConnector[35] = fifoOut[21][3];
              muxOutConnector[36] = fifoOut[22][3];
              muxOutConnector[37] = fifoOut[23][3];
              muxOutConnector[38] = fifoOut[24][3];
              muxOutConnector[39] = fifoOut[25][3];
              muxOutConnector[40] = fifoOut[0][2];
              muxOutConnector[41] = fifoOut[1][2];
              muxOutConnector[42] = fifoOut[2][2];
              muxOutConnector[43] = fifoOut[3][2];
              muxOutConnector[44] = fifoOut[4][2];
              muxOutConnector[45] = fifoOut[5][2];
              muxOutConnector[46] = fifoOut[6][2];
              muxOutConnector[47] = fifoOut[7][2];
              muxOutConnector[48] = fifoOut[8][2];
              muxOutConnector[49] = fifoOut[9][2];
              muxOutConnector[50] = fifoOut[10][2];
              muxOutConnector[51] = fifoOut[11][2];
       end
       11: begin
              muxOutConnector[0] = fifoOut[39][1];
              muxOutConnector[1] = fifoOut[40][1];
              muxOutConnector[2] = fifoOut[41][1];
              muxOutConnector[3] = fifoOut[42][1];
              muxOutConnector[4] = fifoOut[43][1];
              muxOutConnector[5] = fifoOut[44][1];
              muxOutConnector[6] = fifoOut[45][1];
              muxOutConnector[7] = fifoOut[46][1];
              muxOutConnector[8] = fifoOut[47][1];
              muxOutConnector[9] = fifoOut[48][1];
              muxOutConnector[10] = fifoOut[49][1];
              muxOutConnector[11] = fifoOut[50][1];
              muxOutConnector[12] = fifoOut[51][1];
              muxOutConnector[13] = fifoOut[26][0];
              muxOutConnector[14] = fifoOut[27][0];
              muxOutConnector[15] = fifoOut[28][0];
              muxOutConnector[16] = fifoOut[29][0];
              muxOutConnector[17] = fifoOut[30][0];
              muxOutConnector[18] = fifoOut[31][0];
              muxOutConnector[19] = fifoOut[32][0];
              muxOutConnector[20] = fifoOut[33][0];
              muxOutConnector[21] = fifoOut[34][0];
              muxOutConnector[22] = fifoOut[35][0];
              muxOutConnector[23] = fifoOut[36][0];
              muxOutConnector[24] = fifoOut[37][0];
              muxOutConnector[25] = fifoOut[38][0];
              muxOutConnector[26] = fifoOut[12][3];
              muxOutConnector[27] = fifoOut[26][10];
              muxOutConnector[28] = fifoOut[27][10];
              muxOutConnector[29] = fifoOut[28][10];
              muxOutConnector[30] = fifoOut[29][10];
              muxOutConnector[31] = fifoOut[30][10];
              muxOutConnector[32] = fifoOut[31][10];
              muxOutConnector[33] = fifoOut[32][10];
              muxOutConnector[34] = fifoOut[33][10];
              muxOutConnector[35] = fifoOut[34][10];
              muxOutConnector[36] = fifoOut[35][10];
              muxOutConnector[37] = fifoOut[36][10];
              muxOutConnector[38] = fifoOut[37][10];
              muxOutConnector[39] = fifoOut[38][10];
              muxOutConnector[40] = fifoOut[39][10];
              muxOutConnector[41] = fifoOut[40][10];
              muxOutConnector[42] = fifoOut[41][10];
              muxOutConnector[43] = fifoOut[42][10];
              muxOutConnector[44] = fifoOut[43][10];
              muxOutConnector[45] = fifoOut[44][10];
              muxOutConnector[46] = fifoOut[45][10];
              muxOutConnector[47] = fifoOut[46][10];
              muxOutConnector[48] = fifoOut[47][10];
              muxOutConnector[49] = fifoOut[48][10];
              muxOutConnector[50] = fifoOut[49][10];
              muxOutConnector[51] = fifoOut[50][10];
       end
       12: begin
              muxOutConnector[0] = fifoOut[39][1];
              muxOutConnector[1] = fifoOut[40][1];
              muxOutConnector[2] = fifoOut[41][1];
              muxOutConnector[3] = fifoOut[42][1];
              muxOutConnector[4] = fifoOut[43][1];
              muxOutConnector[5] = fifoOut[44][1];
              muxOutConnector[6] = fifoOut[45][1];
              muxOutConnector[7] = fifoOut[46][1];
              muxOutConnector[8] = fifoOut[47][1];
              muxOutConnector[9] = fifoOut[48][1];
              muxOutConnector[10] = fifoOut[49][1];
              muxOutConnector[11] = fifoOut[50][1];
              muxOutConnector[12] = fifoOut[51][1];
              muxOutConnector[13] = fifoOut[26][0];
              muxOutConnector[14] = fifoOut[27][0];
              muxOutConnector[15] = fifoOut[28][0];
              muxOutConnector[16] = fifoOut[29][0];
              muxOutConnector[17] = fifoOut[30][0];
              muxOutConnector[18] = fifoOut[31][0];
              muxOutConnector[19] = fifoOut[32][0];
              muxOutConnector[20] = fifoOut[33][0];
              muxOutConnector[21] = fifoOut[34][0];
              muxOutConnector[22] = fifoOut[35][0];
              muxOutConnector[23] = fifoOut[36][0];
              muxOutConnector[24] = fifoOut[37][0];
              muxOutConnector[25] = fifoOut[38][0];
              muxOutConnector[26] = fifoOut[51][11];
              muxOutConnector[27] = fifoOut[26][10];
              muxOutConnector[28] = fifoOut[27][10];
              muxOutConnector[29] = fifoOut[28][10];
              muxOutConnector[30] = fifoOut[29][10];
              muxOutConnector[31] = fifoOut[30][10];
              muxOutConnector[32] = fifoOut[31][10];
              muxOutConnector[33] = fifoOut[32][10];
              muxOutConnector[34] = fifoOut[33][10];
              muxOutConnector[35] = fifoOut[34][10];
              muxOutConnector[36] = fifoOut[35][10];
              muxOutConnector[37] = fifoOut[36][10];
              muxOutConnector[38] = fifoOut[37][10];
              muxOutConnector[39] = fifoOut[38][10];
              muxOutConnector[40] = fifoOut[39][10];
              muxOutConnector[41] = fifoOut[40][10];
              muxOutConnector[42] = fifoOut[41][10];
              muxOutConnector[43] = fifoOut[42][10];
              muxOutConnector[44] = fifoOut[43][10];
              muxOutConnector[45] = fifoOut[44][10];
              muxOutConnector[46] = fifoOut[45][10];
              muxOutConnector[47] = fifoOut[46][10];
              muxOutConnector[48] = fifoOut[47][10];
              muxOutConnector[49] = fifoOut[48][10];
              muxOutConnector[50] = fifoOut[49][10];
              muxOutConnector[51] = fifoOut[50][10];
       end
       13: begin
              muxOutConnector[0] = fifoOut[39][1];
              muxOutConnector[1] = fifoOut[40][1];
              muxOutConnector[2] = fifoOut[41][1];
              muxOutConnector[3] = fifoOut[42][1];
              muxOutConnector[4] = fifoOut[43][1];
              muxOutConnector[5] = fifoOut[44][1];
              muxOutConnector[6] = fifoOut[45][1];
              muxOutConnector[7] = fifoOut[46][1];
              muxOutConnector[8] = fifoOut[47][1];
              muxOutConnector[9] = fifoOut[48][1];
              muxOutConnector[10] = fifoOut[49][1];
              muxOutConnector[11] = fifoOut[50][1];
              muxOutConnector[12] = fifoOut[51][1];
              muxOutConnector[13] = fifoOut[26][0];
              muxOutConnector[14] = fifoOut[27][0];
              muxOutConnector[15] = fifoOut[28][0];
              muxOutConnector[16] = fifoOut[29][0];
              muxOutConnector[17] = fifoOut[0][12];
              muxOutConnector[18] = fifoOut[1][12];
              muxOutConnector[19] = fifoOut[2][12];
              muxOutConnector[20] = fifoOut[3][12];
              muxOutConnector[21] = fifoOut[4][12];
              muxOutConnector[22] = fifoOut[5][12];
              muxOutConnector[23] = fifoOut[6][12];
              muxOutConnector[24] = fifoOut[7][12];
              muxOutConnector[25] = fifoOut[8][12];
              muxOutConnector[26] = fifoOut[51][11];
              muxOutConnector[27] = fifoOut[26][10];
              muxOutConnector[28] = fifoOut[27][10];
              muxOutConnector[29] = fifoOut[28][10];
              muxOutConnector[30] = fifoOut[29][10];
              muxOutConnector[31] = fifoOut[30][10];
              muxOutConnector[32] = fifoOut[31][10];
              muxOutConnector[33] = fifoOut[32][10];
              muxOutConnector[34] = fifoOut[33][10];
              muxOutConnector[35] = fifoOut[34][10];
              muxOutConnector[36] = fifoOut[35][10];
              muxOutConnector[37] = fifoOut[36][10];
              muxOutConnector[38] = fifoOut[37][10];
              muxOutConnector[39] = fifoOut[38][10];
              muxOutConnector[40] = fifoOut[39][10];
              muxOutConnector[41] = fifoOut[40][10];
              muxOutConnector[42] = fifoOut[41][10];
              muxOutConnector[43] = fifoOut[42][10];
              muxOutConnector[44] = fifoOut[43][10];
              muxOutConnector[45] = fifoOut[44][10];
              muxOutConnector[46] = fifoOut[45][10];
              muxOutConnector[47] = fifoOut[46][10];
              muxOutConnector[48] = fifoOut[47][10];
              muxOutConnector[49] = fifoOut[48][10];
              muxOutConnector[50] = fifoOut[49][10];
              muxOutConnector[51] = fifoOut[50][10];
       end
       14: begin
              muxOutConnector[0] = fifoOut[39][1];
              muxOutConnector[1] = fifoOut[40][1];
              muxOutConnector[2] = fifoOut[41][1];
              muxOutConnector[3] = fifoOut[42][1];
              muxOutConnector[4] = fifoOut[13][0];
              muxOutConnector[5] = fifoOut[14][0];
              muxOutConnector[6] = fifoOut[15][0];
              muxOutConnector[7] = fifoOut[16][0];
              muxOutConnector[8] = fifoOut[17][0];
              muxOutConnector[9] = fifoOut[18][0];
              muxOutConnector[10] = fifoOut[19][0];
              muxOutConnector[11] = fifoOut[20][0];
              muxOutConnector[12] = fifoOut[21][0];
              muxOutConnector[13] = fifoOut[22][0];
              muxOutConnector[14] = fifoOut[23][0];
              muxOutConnector[15] = fifoOut[24][0];
              muxOutConnector[16] = fifoOut[25][0];
              muxOutConnector[17] = fifoOut[0][12];
              muxOutConnector[18] = fifoOut[1][12];
              muxOutConnector[19] = fifoOut[2][12];
              muxOutConnector[20] = fifoOut[3][12];
              muxOutConnector[21] = fifoOut[4][12];
              muxOutConnector[22] = fifoOut[5][12];
              muxOutConnector[23] = fifoOut[6][12];
              muxOutConnector[24] = fifoOut[7][12];
              muxOutConnector[25] = fifoOut[8][12];
              muxOutConnector[26] = fifoOut[51][11];
              muxOutConnector[27] = fifoOut[26][10];
              muxOutConnector[28] = fifoOut[27][10];
              muxOutConnector[29] = fifoOut[28][10];
              muxOutConnector[30] = fifoOut[29][10];
              muxOutConnector[31] = fifoOut[30][10];
              muxOutConnector[32] = fifoOut[31][10];
              muxOutConnector[33] = fifoOut[32][10];
              muxOutConnector[34] = fifoOut[33][10];
              muxOutConnector[35] = fifoOut[34][10];
              muxOutConnector[36] = fifoOut[35][10];
              muxOutConnector[37] = fifoOut[36][10];
              muxOutConnector[38] = fifoOut[37][10];
              muxOutConnector[39] = fifoOut[38][10];
              muxOutConnector[40] = fifoOut[39][10];
              muxOutConnector[41] = fifoOut[40][10];
              muxOutConnector[42] = fifoOut[41][10];
              muxOutConnector[43] = fifoOut[42][10];
              muxOutConnector[44] = fifoOut[43][10];
              muxOutConnector[45] = fifoOut[44][10];
              muxOutConnector[46] = fifoOut[45][10];
              muxOutConnector[47] = fifoOut[46][10];
              muxOutConnector[48] = fifoOut[47][10];
              muxOutConnector[49] = fifoOut[48][10];
              muxOutConnector[50] = fifoOut[49][10];
              muxOutConnector[51] = fifoOut[50][10];
       end
       15: begin
              muxOutConnector[0] = fifoOut[9][0];
              muxOutConnector[1] = fifoOut[10][0];
              muxOutConnector[2] = fifoOut[11][0];
              muxOutConnector[3] = fifoOut[12][0];
              muxOutConnector[4] = fifoOut[13][0];
              muxOutConnector[5] = fifoOut[14][0];
              muxOutConnector[6] = fifoOut[15][0];
              muxOutConnector[7] = fifoOut[16][0];
              muxOutConnector[8] = fifoOut[17][0];
              muxOutConnector[9] = fifoOut[18][0];
              muxOutConnector[10] = fifoOut[19][0];
              muxOutConnector[11] = fifoOut[20][0];
              muxOutConnector[12] = fifoOut[21][0];
              muxOutConnector[13] = fifoOut[22][0];
              muxOutConnector[14] = fifoOut[23][0];
              muxOutConnector[15] = fifoOut[24][0];
              muxOutConnector[16] = fifoOut[25][0];
              muxOutConnector[17] = fifoOut[0][12];
              muxOutConnector[18] = fifoOut[1][12];
              muxOutConnector[19] = fifoOut[2][12];
              muxOutConnector[20] = fifoOut[3][12];
              muxOutConnector[21] = fifoOut[4][12];
              muxOutConnector[22] = fifoOut[5][12];
              muxOutConnector[23] = fifoOut[6][12];
              muxOutConnector[24] = fifoOut[7][12];
              muxOutConnector[25] = fifoOut[8][12];
              muxOutConnector[26] = fifoOut[51][11];
              muxOutConnector[27] = fifoOut[26][10];
              muxOutConnector[28] = fifoOut[27][10];
              muxOutConnector[29] = fifoOut[28][10];
              muxOutConnector[30] = fifoOut[29][10];
              muxOutConnector[31] = fifoOut[30][10];
              muxOutConnector[32] = fifoOut[31][10];
              muxOutConnector[33] = fifoOut[32][10];
              muxOutConnector[34] = fifoOut[33][10];
              muxOutConnector[35] = fifoOut[34][10];
              muxOutConnector[36] = fifoOut[35][10];
              muxOutConnector[37] = fifoOut[36][10];
              muxOutConnector[38] = fifoOut[37][10];
              muxOutConnector[39] = fifoOut[38][10];
              muxOutConnector[40] = fifoOut[39][10];
              muxOutConnector[41] = fifoOut[40][10];
              muxOutConnector[42] = fifoOut[41][10];
              muxOutConnector[43] = fifoOut[42][10];
              muxOutConnector[44] = fifoOut[43][10];
              muxOutConnector[45] = fifoOut[44][10];
              muxOutConnector[46] = fifoOut[45][10];
              muxOutConnector[47] = fifoOut[46][10];
              muxOutConnector[48] = fifoOut[47][10];
              muxOutConnector[49] = fifoOut[48][10];
              muxOutConnector[50] = fifoOut[49][10];
              muxOutConnector[51] = fifoOut[50][10];
       end
       16: begin
              muxOutConnector[0] = fifoOut[9][0];
              muxOutConnector[1] = fifoOut[10][0];
              muxOutConnector[2] = fifoOut[11][0];
              muxOutConnector[3] = fifoOut[12][0];
              muxOutConnector[4] = fifoOut[13][0];
              muxOutConnector[5] = fifoOut[14][0];
              muxOutConnector[6] = fifoOut[15][0];
              muxOutConnector[7] = fifoOut[16][0];
              muxOutConnector[8] = fifoOut[17][0];
              muxOutConnector[9] = fifoOut[18][0];
              muxOutConnector[10] = fifoOut[19][0];
              muxOutConnector[11] = fifoOut[20][0];
              muxOutConnector[12] = fifoOut[21][0];
              muxOutConnector[13] = fifoOut[22][0];
              muxOutConnector[14] = fifoOut[23][0];
              muxOutConnector[15] = fifoOut[24][0];
              muxOutConnector[16] = fifoOut[25][0];
              muxOutConnector[17] = fifoOut[0][12];
              muxOutConnector[18] = fifoOut[1][12];
              muxOutConnector[19] = fifoOut[2][12];
              muxOutConnector[20] = fifoOut[3][12];
              muxOutConnector[21] = fifoOut[4][12];
              muxOutConnector[22] = fifoOut[5][12];
              muxOutConnector[23] = fifoOut[6][12];
              muxOutConnector[24] = fifoOut[7][12];
              muxOutConnector[25] = fifoOut[8][12];
              muxOutConnector[26] = fifoOut[51][11];
              muxOutConnector[27] = fifoOut[26][10];
              muxOutConnector[28] = fifoOut[27][10];
              muxOutConnector[29] = fifoOut[28][10];
              muxOutConnector[30] = fifoOut[29][10];
              muxOutConnector[31] = fifoOut[30][10];
              muxOutConnector[32] = fifoOut[31][10];
              muxOutConnector[33] = fifoOut[32][10];
              muxOutConnector[34] = fifoOut[33][10];
              muxOutConnector[35] = fifoOut[34][10];
              muxOutConnector[36] = fifoOut[35][10];
              muxOutConnector[37] = fifoOut[36][10];
              muxOutConnector[38] = fifoOut[37][10];
              muxOutConnector[39] = fifoOut[38][10];
              muxOutConnector[40] = fifoOut[39][10];
              muxOutConnector[41] = fifoOut[40][10];
              muxOutConnector[42] = fifoOut[41][10];
              muxOutConnector[43] = fifoOut[42][10];
              muxOutConnector[44] = fifoOut[43][10];
              muxOutConnector[45] = fifoOut[44][10];
              muxOutConnector[46] = fifoOut[45][10];
              muxOutConnector[47] = fifoOut[46][10];
              muxOutConnector[48] = fifoOut[47][10];
              muxOutConnector[49] = fifoOut[48][10];
              muxOutConnector[50] = fifoOut[49][10];
              muxOutConnector[51] = fifoOut[50][10];
       end
       17: begin
              muxOutConnector[0] = fifoOut[9][0];
              muxOutConnector[1] = fifoOut[10][0];
              muxOutConnector[2] = fifoOut[11][0];
              muxOutConnector[3] = fifoOut[12][0];
              muxOutConnector[4] = fifoOut[13][0];
              muxOutConnector[5] = fifoOut[14][0];
              muxOutConnector[6] = fifoOut[15][0];
              muxOutConnector[7] = fifoOut[16][0];
              muxOutConnector[8] = fifoOut[17][0];
              muxOutConnector[9] = fifoOut[18][0];
              muxOutConnector[10] = fifoOut[19][0];
              muxOutConnector[11] = fifoOut[20][0];
              muxOutConnector[12] = fifoOut[21][0];
              muxOutConnector[13] = fifoOut[22][0];
              muxOutConnector[14] = fifoOut[23][0];
              muxOutConnector[15] = fifoOut[24][0];
              muxOutConnector[16] = fifoOut[25][0];
              muxOutConnector[17] = fifoOut[0][12];
              muxOutConnector[18] = fifoOut[1][12];
              muxOutConnector[19] = fifoOut[2][12];
              muxOutConnector[20] = fifoOut[3][12];
              muxOutConnector[21] = fifoOut[4][12];
              muxOutConnector[22] = fifoOut[5][12];
              muxOutConnector[23] = fifoOut[6][12];
              muxOutConnector[24] = fifoOut[7][12];
              muxOutConnector[25] = fifoOut[8][12];
              muxOutConnector[26] = fifoOut[51][11];
              muxOutConnector[27] = fifoOut[26][10];
              muxOutConnector[28] = fifoOut[27][10];
              muxOutConnector[29] = fifoOut[28][10];
              muxOutConnector[30] = fifoOut[29][10];
              muxOutConnector[31] = fifoOut[30][10];
              muxOutConnector[32] = fifoOut[31][10];
              muxOutConnector[33] = fifoOut[32][10];
              muxOutConnector[34] = fifoOut[33][10];
              muxOutConnector[35] = fifoOut[34][10];
              muxOutConnector[36] = fifoOut[35][10];
              muxOutConnector[37] = fifoOut[36][10];
              muxOutConnector[38] = fifoOut[37][10];
              muxOutConnector[39] = fifoOut[38][10];
              muxOutConnector[40] = fifoOut[39][10];
              muxOutConnector[41] = fifoOut[40][10];
              muxOutConnector[42] = fifoOut[41][10];
              muxOutConnector[43] = fifoOut[42][10];
              muxOutConnector[44] = fifoOut[43][10];
              muxOutConnector[45] = fifoOut[44][10];
              muxOutConnector[46] = fifoOut[45][10];
              muxOutConnector[47] = fifoOut[46][10];
              muxOutConnector[48] = fifoOut[47][10];
              muxOutConnector[49] = fifoOut[48][10];
              muxOutConnector[50] = fifoOut[49][10];
              muxOutConnector[51] = fifoOut[50][10];
       end
       18: begin
              muxOutConnector[0] = fifoOut[9][0];
              muxOutConnector[1] = fifoOut[10][0];
              muxOutConnector[2] = fifoOut[11][0];
              muxOutConnector[3] = fifoOut[12][0];
              muxOutConnector[4] = fifoOut[13][0];
              muxOutConnector[5] = fifoOut[14][0];
              muxOutConnector[6] = fifoOut[15][0];
              muxOutConnector[7] = fifoOut[16][0];
              muxOutConnector[8] = fifoOut[17][0];
              muxOutConnector[9] = fifoOut[18][0];
              muxOutConnector[10] = fifoOut[19][0];
              muxOutConnector[11] = fifoOut[20][0];
              muxOutConnector[12] = fifoOut[21][0];
              muxOutConnector[13] = fifoOut[22][0];
              muxOutConnector[14] = fifoOut[23][0];
              muxOutConnector[15] = fifoOut[24][0];
              muxOutConnector[16] = fifoOut[25][0];
              muxOutConnector[17] = fifoOut[0][12];
              muxOutConnector[18] = fifoOut[1][12];
              muxOutConnector[19] = fifoOut[2][12];
              muxOutConnector[20] = fifoOut[3][12];
              muxOutConnector[21] = fifoOut[4][12];
              muxOutConnector[22] = fifoOut[5][12];
              muxOutConnector[23] = fifoOut[6][12];
              muxOutConnector[24] = fifoOut[7][12];
              muxOutConnector[25] = fifoOut[8][12];
              muxOutConnector[26] = fifoOut[51][11];
              muxOutConnector[27] = fifoOut[26][10];
              muxOutConnector[28] = fifoOut[27][10];
              muxOutConnector[29] = fifoOut[28][10];
              muxOutConnector[30] = fifoOut[29][10];
              muxOutConnector[31] = fifoOut[30][10];
              muxOutConnector[32] = fifoOut[31][10];
              muxOutConnector[33] = fifoOut[32][10];
              muxOutConnector[34] = fifoOut[33][10];
              muxOutConnector[35] = fifoOut[34][10];
              muxOutConnector[36] = fifoOut[35][10];
              muxOutConnector[37] = fifoOut[36][10];
              muxOutConnector[38] = fifoOut[37][10];
              muxOutConnector[39] = fifoOut[38][10];
              muxOutConnector[40] = fifoOut[39][10];
              muxOutConnector[41] = fifoOut[40][10];
              muxOutConnector[42] = fifoOut[41][10];
              muxOutConnector[43] = fifoOut[42][10];
              muxOutConnector[44] = fifoOut[43][10];
              muxOutConnector[45] = fifoOut[44][10];
              muxOutConnector[46] = fifoOut[45][10];
              muxOutConnector[47] = fifoOut[46][10];
              muxOutConnector[48] = fifoOut[47][10];
              muxOutConnector[49] = fifoOut[48][10];
              muxOutConnector[50] = fifoOut[49][10];
              muxOutConnector[51] = fifoOut[50][10];
       end
       19: begin
              muxOutConnector[0] = fifoOut[9][0];
              muxOutConnector[1] = fifoOut[10][0];
              muxOutConnector[2] = fifoOut[11][0];
              muxOutConnector[3] = fifoOut[12][0];
              muxOutConnector[4] = fifoOut[13][0];
              muxOutConnector[5] = fifoOut[14][0];
              muxOutConnector[6] = fifoOut[15][0];
              muxOutConnector[7] = fifoOut[16][0];
              muxOutConnector[8] = fifoOut[17][0];
              muxOutConnector[9] = fifoOut[18][0];
              muxOutConnector[10] = fifoOut[19][0];
              muxOutConnector[11] = fifoOut[20][0];
              muxOutConnector[12] = fifoOut[21][0];
              muxOutConnector[13] = fifoOut[22][0];
              muxOutConnector[14] = fifoOut[23][0];
              muxOutConnector[15] = fifoOut[24][0];
              muxOutConnector[16] = fifoOut[25][0];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[51][11];
              muxOutConnector[27] = fifoOut[26][10];
              muxOutConnector[28] = fifoOut[27][10];
              muxOutConnector[29] = fifoOut[28][10];
              muxOutConnector[30] = fifoOut[29][10];
              muxOutConnector[31] = fifoOut[30][10];
              muxOutConnector[32] = fifoOut[31][10];
              muxOutConnector[33] = fifoOut[32][10];
              muxOutConnector[34] = fifoOut[33][10];
              muxOutConnector[35] = fifoOut[34][10];
              muxOutConnector[36] = fifoOut[35][10];
              muxOutConnector[37] = fifoOut[36][10];
              muxOutConnector[38] = fifoOut[37][10];
              muxOutConnector[39] = fifoOut[38][10];
              muxOutConnector[40] = fifoOut[39][10];
              muxOutConnector[41] = fifoOut[40][10];
              muxOutConnector[42] = fifoOut[41][10];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
