`timescale 1ns / 1ps
module Dmem_circ8_scripted(
		 muxOut,
		 dMemIn,
		 wr_en,
		 reaccessAddress,
		 reaccess_lyr,
		 rd_en, clk, rst 
 );
parameter r = 52;
parameter c = 12;
parameter w = 6;
parameter ADDRESSWIDTH = 5;

parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 
output wire [r*w -1 : 0]muxOut;// r numbers of w bits
input [r*w-1:0]dMemIn;
input wr_en;
input [ADDRESSWIDTH-1:0]reaccessAddress;
input reaccess_lyr;
input rd_en;
input clk,rst;

wire [(ADDRESSWIDTH+1)-1:0]case_sel;//{layer,address}
wire [w-1:0]dMemInDummy[r-1:0];
reg [w-1:0]muxOutWire[r-1:0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<r;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutWire[k];
        assign dMemInDummy[k] = dMemIn[ (k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always @(posedge clk) begin
    if (rst) begin
         for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] = 0;
           end
        end
    end
    else begin
    if(wr_en) begin
        // Set (i,j)th value = (i,j-1)th value
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Load Inputs
        for(i = r-1; i > -1; i=i-1) begin
            fifoOut[i][0] <= dMemInDummy[i]; 
        end
    end
    else begin 
        // Set (i,j)th value = (i,j)th value
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <= fifoOut[i][j];
            end
        end
    end
    end
end

assign case_sel = rd_en ? {reaccess_lyr,reaccessAddress} : {1'd1,READDISABLEDCASE};

always@(*) begin
    case(case_sel)

		 {1'd0, 5'd0} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd1} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd2} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd3} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd4} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd5} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd6} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd7} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 4 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 4 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 4 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 4 ]; 
		 end
		 {1'd0, 5'd8} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 5 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 5 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 5 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 5 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 5 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 5 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 5 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 5 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 5 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 5 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 5 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 5 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 5 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 5 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 5 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 5 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 5 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 5 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 5 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 5 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 5 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 5 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 4 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 4 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 4 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 4 ]; 
		 end
		 {1'd0, 5'd9} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 5 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 5 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 5 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 5 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 5 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 5 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 5 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 5 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 5 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 5 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 5 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 5 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 5 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 5 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 5 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 5 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 5 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 5 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 5 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 5 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 5 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 5 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 4 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 4 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 4 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 4 ]; 
		 end
		 {1'd0, 5'd10} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 5 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 5 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 5 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 5 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 5 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 5 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 5 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 5 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 5 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 5 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 5 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 5 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 5 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 5 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 5 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 5 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 5 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 5 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 5 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 5 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 5 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 5 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 4 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 4 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 4 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 4 ]; 
		 end
		 {1'd0, 5'd11} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 8 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 8 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 8 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 8 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 8 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 5 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 5 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 5 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 5 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 5 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 5 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 5 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 5 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 5 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 5 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 5 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 5 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 5 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 5 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 5 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 5 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 5 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 5 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 5 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 5 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 5 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 5 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 4 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 4 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 4 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 4 ]; 
		 end
		 {1'd0, 5'd12} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 9 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 9 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 9 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 9 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 9 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 9 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 9 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 9 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 9 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 9 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 9 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 9 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 9 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 9 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 9 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 9 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 9 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 9 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 9 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 9 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 9 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 8 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 8 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 8 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 8 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 8 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 5 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 5 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 5 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 5 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 5 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 5 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 5 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 5 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 5 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 5 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 5 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 5 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 5 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 5 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 5 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 5 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 5 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 5 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 5 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 5 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 5 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 5 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 4 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 4 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 4 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 4 ]; 
		 end
		 {1'd0, 5'd13} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 9 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 9 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 9 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 9 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 9 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 9 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 9 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 9 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 9 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 9 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 9 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 9 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 9 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 9 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 9 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 9 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 9 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 9 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 9 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 9 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 9 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 8 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 8 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 8 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 8 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 8 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 5 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 5 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 5 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 5 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 5 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 5 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 5 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 5 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 5 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 5 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 5 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 5 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 5 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 5 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 5 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 5 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 5 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 5 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 5 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 5 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 5 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 5 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 4 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 4 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 4 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 4 ]; 
		 end
		 {1'd0, 5'd14} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 9 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 9 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 9 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 9 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 9 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 9 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 9 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 9 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 9 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 9 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 9 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 9 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 9 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 9 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 9 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 9 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 9 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 9 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 9 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 9 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 9 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 8 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 8 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 8 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 8 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 8 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 5 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 5 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 5 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 5 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 5 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 5 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 5 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 5 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 5 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 5 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 5 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 5 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 5 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 5 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 5 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 5 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 5 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 5 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 5 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 5 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 5 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 5 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 4 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 4 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 4 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 4 ]; 
		 end
		 {1'd0, 5'd15} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 9 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 9 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 9 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 9 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 9 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 9 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 9 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 9 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 9 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 9 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 9 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 9 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 9 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 9 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 9 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 9 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 9 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 9 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 9 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 9 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 9 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 8 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 8 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 8 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 8 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 8 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 5 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 5 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 5 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 5 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 5 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 5 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 5 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 5 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 5 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 5 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 5 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 5 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 5 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 5 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 5 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 5 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 5 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 5 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 5 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 5 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 5 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 5 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 4 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 4 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 4 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 4 ]; 
		 end
		 {1'd0, 5'd16} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 9 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 9 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 9 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 9 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 9 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 9 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 9 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 9 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 9 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 9 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 9 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 9 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 9 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 9 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 9 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 9 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 9 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 9 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 9 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 9 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 9 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 8 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 8 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 8 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 8 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 8 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 5 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 5 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 5 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 5 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 5 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 5 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 5 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 5 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 5 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 5 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 5 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 5 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 5 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 5 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 5 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 5 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 5 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 5 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 5 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 5 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 5 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 5 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 4 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 4 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 4 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 4 ]; 
		 end
		 {1'd0, 5'd17} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 9 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 9 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 9 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 9 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 9 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 9 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 9 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 9 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 9 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 9 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 9 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 9 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 9 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 9 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 9 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 9 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 9 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 9 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 9 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 9 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 9 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 8 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 8 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 8 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 8 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 8 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 5 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 5 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 5 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 5 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 5 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 5 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 5 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 5 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 5 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 5 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 5 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 5 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 5 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 5 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 5 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 5 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 5 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 5 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 5 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 5 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 5 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 5 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 4 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 4 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 4 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 4 ]; 
		 end
		 {1'd0, 5'd18} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 9 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 9 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 9 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 9 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 9 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 9 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 9 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 9 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 9 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 9 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 9 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 9 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 9 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 9 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 9 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 9 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 9 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 9 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 9 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 9 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 9 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 8 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 8 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 8 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 8 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 8 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 5 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 5 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 5 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 5 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 5 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 5 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 5 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 5 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 5 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 5 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 5 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 5 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 5 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 5 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 5 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 5 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 5 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 5 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 5 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 5 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 5 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 5 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 4 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 4 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 4 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 4 ]; 
		 end
		 {1'd0, 5'd19} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 9 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 9 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 9 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 9 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 9 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 9 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 9 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 9 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 9 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 9 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 9 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 9 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 9 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 9 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 9 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 9 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 9 ]; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 5 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 5 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 5 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 5 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 5 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 5 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 5 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 5 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 5 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 5 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 5 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 5 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 5 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 5 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 5 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 5 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 5 ]; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd0} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd1} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd2} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd3} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd4} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd5} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd6} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 32 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd7} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 32 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd8} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 32 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd9} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 32 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd10} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 32 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd11} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 32 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd12} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 32 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd13} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 32 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = fifoOut[ 0 ][ 10 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 1 ][ 10 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 2 ][ 10 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 3 ][ 10 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 4 ][ 10 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 5 ][ 10 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 6 ][ 10 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 7 ][ 10 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 8 ][ 10 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 9 ][ 10 ]; 
		 end
		 {1'd1, 5'd14} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 32 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 10 ][ 11 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 11 ][ 11 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 12 ][ 11 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 13 ][ 11 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 14 ][ 11 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 15 ][ 11 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 16 ][ 11 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 17 ][ 11 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 18 ][ 11 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 19 ][ 11 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 20 ][ 11 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 21 ][ 11 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 22 ][ 11 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 23 ][ 11 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 24 ][ 11 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 25 ][ 11 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 0 ][ 10 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 1 ][ 10 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 2 ][ 10 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 3 ][ 10 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 4 ][ 10 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 5 ][ 10 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 6 ][ 10 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 7 ][ 10 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 8 ][ 10 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 9 ][ 10 ]; 
		 end
		 {1'd1, 5'd15} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 32 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 10 ][ 11 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 11 ][ 11 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 12 ][ 11 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 13 ][ 11 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 14 ][ 11 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 15 ][ 11 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 16 ][ 11 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 17 ][ 11 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 18 ][ 11 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 19 ][ 11 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 20 ][ 11 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 21 ][ 11 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 22 ][ 11 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 23 ][ 11 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 24 ][ 11 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 25 ][ 11 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 0 ][ 10 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 1 ][ 10 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 2 ][ 10 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 3 ][ 10 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 4 ][ 10 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 5 ][ 10 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 6 ][ 10 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 7 ][ 10 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 8 ][ 10 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 9 ][ 10 ]; 
		 end
		 {1'd1, 5'd16} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 32 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 10 ][ 11 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 11 ][ 11 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 12 ][ 11 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 13 ][ 11 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 14 ][ 11 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 15 ][ 11 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 16 ][ 11 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 17 ][ 11 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 18 ][ 11 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 19 ][ 11 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 20 ][ 11 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 21 ][ 11 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 22 ][ 11 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 23 ][ 11 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 24 ][ 11 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 25 ][ 11 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 0 ][ 10 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 1 ][ 10 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 2 ][ 10 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 3 ][ 10 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 4 ][ 10 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 5 ][ 10 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 6 ][ 10 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 7 ][ 10 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 8 ][ 10 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 9 ][ 10 ]; 
		 end
		 {1'd1, 5'd17} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 32 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 10 ][ 11 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 11 ][ 11 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 12 ][ 11 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 13 ][ 11 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 14 ][ 11 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 15 ][ 11 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 16 ][ 11 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 17 ][ 11 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 18 ][ 11 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 19 ][ 11 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 20 ][ 11 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 21 ][ 11 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 22 ][ 11 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 23 ][ 11 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 24 ][ 11 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 25 ][ 11 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 0 ][ 10 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 1 ][ 10 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 2 ][ 10 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 3 ][ 10 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 4 ][ 10 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 5 ][ 10 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 6 ][ 10 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 7 ][ 10 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 8 ][ 10 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 9 ][ 10 ]; 
		 end
		 {1'd1, 5'd18} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 32 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 42 ][ 3 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 43 ][ 3 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 44 ][ 3 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 45 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 46 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 47 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 48 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 49 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 50 ][ 3 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 10 ][ 11 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 11 ][ 11 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 12 ][ 11 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 13 ][ 11 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 14 ][ 11 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 15 ][ 11 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 16 ][ 11 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 17 ][ 11 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 18 ][ 11 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 19 ][ 11 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 20 ][ 11 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 21 ][ 11 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 22 ][ 11 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 23 ][ 11 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 24 ][ 11 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 25 ][ 11 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 0 ][ 10 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 1 ][ 10 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 2 ][ 10 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 3 ][ 10 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 4 ][ 10 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 5 ][ 10 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 6 ][ 10 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 7 ][ 10 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 8 ][ 10 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 9 ][ 10 ]; 
		 end
		 {1'd1, 5'd19} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 32 ][ 3 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 33 ][ 3 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 34 ][ 3 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 35 ][ 3 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 36 ][ 3 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 37 ][ 3 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 38 ][ 3 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 39 ][ 3 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 40 ][ 3 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 41 ][ 3 ]; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 10 ][ 11 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 11 ][ 11 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 12 ][ 11 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 13 ][ 11 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 14 ][ 11 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 15 ][ 11 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 16 ][ 11 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 17 ][ 11 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 18 ][ 11 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 19 ][ 11 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 20 ][ 11 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 21 ][ 11 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 22 ][ 11 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 23 ][ 11 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 24 ][ 11 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 25 ][ 11 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 0 ][ 10 ]; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
    default:begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
    end
    endcase
end
endmodule
