`timescale 1ns / 1ps
module LMem0To1_511_circ4_ys_scripted(
        muxOut,
        ly0In,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 16;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

reg   feedback_en;
reg [ w - 1 : 0 ]column_1[ r - 1 : 0 ];
reg chip_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(chip_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= column_1[i];
         end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
  feedback_en=rd_en;
      if(wr_en)begin
        chip_en=wr_en;
      end
      else begin
        chip_en=feedback_en;
      end
   if(feedback_en)begin
      for(i = r-1; i > -1; i=i-1) begin
        column_1[i] = fifoOut[i][c-1];
      end
   end
   else begin
      for(i = r-1; i > -1; i=i-1) begin
        column_1[i] = ly0InConnector[i];
      end
    end
end
always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[7][11];
              muxOutConnector[1] = fifoOut[8][11];
              muxOutConnector[2] = fifoOut[9][11];
              muxOutConnector[3] = fifoOut[10][11];
              muxOutConnector[4] = fifoOut[11][11];
              muxOutConnector[5] = fifoOut[12][11];
              muxOutConnector[6] = fifoOut[13][11];
              muxOutConnector[7] = fifoOut[14][11];
              muxOutConnector[8] = fifoOut[15][11];
              muxOutConnector[9] = fifoOut[16][11];
              muxOutConnector[10] = fifoOut[17][11];
              muxOutConnector[11] = fifoOut[18][11];
              muxOutConnector[12] = fifoOut[19][11];
              muxOutConnector[13] = fifoOut[20][11];
              muxOutConnector[14] = fifoOut[21][11];
              muxOutConnector[15] = fifoOut[22][11];
              muxOutConnector[16] = fifoOut[23][11];
              muxOutConnector[17] = fifoOut[24][11];
              muxOutConnector[18] = fifoOut[25][11];
              muxOutConnector[19] = fifoOut[0][10];
              muxOutConnector[20] = fifoOut[1][10];
              muxOutConnector[21] = fifoOut[2][10];
              muxOutConnector[22] = fifoOut[3][10];
              muxOutConnector[23] = fifoOut[4][10];
              muxOutConnector[24] = fifoOut[5][10];
              muxOutConnector[25] = fifoOut[6][10];
              muxOutConnector[26] = fifoOut[4][3];
              muxOutConnector[27] = fifoOut[5][3];
              muxOutConnector[28] = fifoOut[6][3];
              muxOutConnector[29] = fifoOut[7][3];
              muxOutConnector[30] = fifoOut[8][3];
              muxOutConnector[31] = fifoOut[9][3];
              muxOutConnector[32] = fifoOut[10][3];
              muxOutConnector[33] = fifoOut[11][3];
              muxOutConnector[34] = fifoOut[12][3];
              muxOutConnector[35] = fifoOut[13][3];
              muxOutConnector[36] = fifoOut[14][3];
              muxOutConnector[37] = fifoOut[15][3];
              muxOutConnector[38] = fifoOut[16][3];
              muxOutConnector[39] = fifoOut[17][3];
              muxOutConnector[40] = fifoOut[18][3];
              muxOutConnector[41] = fifoOut[19][3];
              muxOutConnector[42] = fifoOut[20][3];
              muxOutConnector[43] = fifoOut[21][3];
              muxOutConnector[44] = fifoOut[22][3];
              muxOutConnector[45] = fifoOut[23][3];
              muxOutConnector[46] = fifoOut[24][3];
              muxOutConnector[47] = fifoOut[25][3];
              muxOutConnector[48] = fifoOut[0][2];
              muxOutConnector[49] = fifoOut[1][2];
              muxOutConnector[50] = fifoOut[2][2];
              muxOutConnector[51] = fifoOut[3][2];
       end
       1: begin
              muxOutConnector[0] = fifoOut[7][11];
              muxOutConnector[1] = fifoOut[8][11];
              muxOutConnector[2] = fifoOut[9][11];
              muxOutConnector[3] = fifoOut[10][11];
              muxOutConnector[4] = fifoOut[11][11];
              muxOutConnector[5] = fifoOut[12][11];
              muxOutConnector[6] = fifoOut[13][11];
              muxOutConnector[7] = fifoOut[14][11];
              muxOutConnector[8] = fifoOut[15][11];
              muxOutConnector[9] = fifoOut[16][11];
              muxOutConnector[10] = fifoOut[17][11];
              muxOutConnector[11] = fifoOut[18][11];
              muxOutConnector[12] = fifoOut[19][11];
              muxOutConnector[13] = fifoOut[20][11];
              muxOutConnector[14] = fifoOut[21][11];
              muxOutConnector[15] = fifoOut[22][11];
              muxOutConnector[16] = fifoOut[23][11];
              muxOutConnector[17] = fifoOut[24][11];
              muxOutConnector[18] = fifoOut[25][11];
              muxOutConnector[19] = fifoOut[0][10];
              muxOutConnector[20] = fifoOut[1][10];
              muxOutConnector[21] = fifoOut[2][10];
              muxOutConnector[22] = fifoOut[3][10];
              muxOutConnector[23] = fifoOut[4][10];
              muxOutConnector[24] = fifoOut[5][10];
              muxOutConnector[25] = fifoOut[6][10];
              muxOutConnector[26] = fifoOut[4][3];
              muxOutConnector[27] = fifoOut[5][3];
              muxOutConnector[28] = fifoOut[6][3];
              muxOutConnector[29] = fifoOut[7][3];
              muxOutConnector[30] = fifoOut[8][3];
              muxOutConnector[31] = fifoOut[9][3];
              muxOutConnector[32] = fifoOut[10][3];
              muxOutConnector[33] = fifoOut[11][3];
              muxOutConnector[34] = fifoOut[12][3];
              muxOutConnector[35] = fifoOut[13][3];
              muxOutConnector[36] = fifoOut[14][3];
              muxOutConnector[37] = fifoOut[15][3];
              muxOutConnector[38] = fifoOut[16][3];
              muxOutConnector[39] = fifoOut[17][3];
              muxOutConnector[40] = fifoOut[18][3];
              muxOutConnector[41] = fifoOut[19][3];
              muxOutConnector[42] = fifoOut[20][3];
              muxOutConnector[43] = fifoOut[21][3];
              muxOutConnector[44] = fifoOut[22][3];
              muxOutConnector[45] = fifoOut[23][3];
              muxOutConnector[46] = fifoOut[24][3];
              muxOutConnector[47] = fifoOut[25][3];
              muxOutConnector[48] = fifoOut[0][2];
              muxOutConnector[49] = fifoOut[1][2];
              muxOutConnector[50] = fifoOut[2][2];
              muxOutConnector[51] = fifoOut[3][2];
       end
       2: begin
              muxOutConnector[0] = fifoOut[7][11];
              muxOutConnector[1] = fifoOut[8][11];
              muxOutConnector[2] = fifoOut[9][11];
              muxOutConnector[3] = fifoOut[10][11];
              muxOutConnector[4] = fifoOut[11][11];
              muxOutConnector[5] = fifoOut[12][11];
              muxOutConnector[6] = fifoOut[13][11];
              muxOutConnector[7] = fifoOut[14][11];
              muxOutConnector[8] = fifoOut[15][11];
              muxOutConnector[9] = fifoOut[16][11];
              muxOutConnector[10] = fifoOut[17][11];
              muxOutConnector[11] = fifoOut[18][11];
              muxOutConnector[12] = fifoOut[19][11];
              muxOutConnector[13] = fifoOut[20][11];
              muxOutConnector[14] = fifoOut[21][11];
              muxOutConnector[15] = fifoOut[22][11];
              muxOutConnector[16] = fifoOut[23][11];
              muxOutConnector[17] = fifoOut[24][11];
              muxOutConnector[18] = fifoOut[25][11];
              muxOutConnector[19] = fifoOut[0][10];
              muxOutConnector[20] = fifoOut[1][10];
              muxOutConnector[21] = fifoOut[2][10];
              muxOutConnector[22] = fifoOut[3][10];
              muxOutConnector[23] = fifoOut[4][10];
              muxOutConnector[24] = fifoOut[5][10];
              muxOutConnector[25] = fifoOut[6][10];
              muxOutConnector[26] = fifoOut[4][3];
              muxOutConnector[27] = fifoOut[5][3];
              muxOutConnector[28] = fifoOut[6][3];
              muxOutConnector[29] = fifoOut[7][3];
              muxOutConnector[30] = fifoOut[8][3];
              muxOutConnector[31] = fifoOut[9][3];
              muxOutConnector[32] = fifoOut[10][3];
              muxOutConnector[33] = fifoOut[11][3];
              muxOutConnector[34] = fifoOut[12][3];
              muxOutConnector[35] = fifoOut[13][3];
              muxOutConnector[36] = fifoOut[14][3];
              muxOutConnector[37] = fifoOut[15][3];
              muxOutConnector[38] = fifoOut[16][3];
              muxOutConnector[39] = fifoOut[17][3];
              muxOutConnector[40] = fifoOut[18][3];
              muxOutConnector[41] = fifoOut[19][3];
              muxOutConnector[42] = fifoOut[20][3];
              muxOutConnector[43] = fifoOut[21][3];
              muxOutConnector[44] = fifoOut[22][3];
              muxOutConnector[45] = fifoOut[23][3];
              muxOutConnector[46] = fifoOut[24][3];
              muxOutConnector[47] = fifoOut[25][3];
              muxOutConnector[48] = fifoOut[0][2];
              muxOutConnector[49] = fifoOut[1][2];
              muxOutConnector[50] = fifoOut[2][2];
              muxOutConnector[51] = fifoOut[3][2];
       end
       3: begin
              muxOutConnector[0] = fifoOut[7][11];
              muxOutConnector[1] = fifoOut[8][11];
              muxOutConnector[2] = fifoOut[9][11];
              muxOutConnector[3] = fifoOut[10][11];
              muxOutConnector[4] = fifoOut[11][11];
              muxOutConnector[5] = fifoOut[12][11];
              muxOutConnector[6] = fifoOut[13][11];
              muxOutConnector[7] = fifoOut[14][11];
              muxOutConnector[8] = fifoOut[15][11];
              muxOutConnector[9] = fifoOut[16][11];
              muxOutConnector[10] = fifoOut[17][11];
              muxOutConnector[11] = fifoOut[18][11];
              muxOutConnector[12] = fifoOut[19][11];
              muxOutConnector[13] = fifoOut[20][11];
              muxOutConnector[14] = fifoOut[21][11];
              muxOutConnector[15] = fifoOut[22][11];
              muxOutConnector[16] = fifoOut[23][11];
              muxOutConnector[17] = fifoOut[24][11];
              muxOutConnector[18] = fifoOut[25][11];
              muxOutConnector[19] = fifoOut[0][10];
              muxOutConnector[20] = fifoOut[1][10];
              muxOutConnector[21] = fifoOut[2][10];
              muxOutConnector[22] = fifoOut[3][10];
              muxOutConnector[23] = fifoOut[4][10];
              muxOutConnector[24] = fifoOut[5][10];
              muxOutConnector[25] = fifoOut[6][10];
              muxOutConnector[26] = fifoOut[4][3];
              muxOutConnector[27] = fifoOut[5][3];
              muxOutConnector[28] = fifoOut[6][3];
              muxOutConnector[29] = fifoOut[7][3];
              muxOutConnector[30] = fifoOut[8][3];
              muxOutConnector[31] = fifoOut[9][3];
              muxOutConnector[32] = fifoOut[10][3];
              muxOutConnector[33] = fifoOut[11][3];
              muxOutConnector[34] = fifoOut[12][3];
              muxOutConnector[35] = fifoOut[13][3];
              muxOutConnector[36] = fifoOut[14][3];
              muxOutConnector[37] = fifoOut[15][3];
              muxOutConnector[38] = fifoOut[16][3];
              muxOutConnector[39] = fifoOut[41][2];
              muxOutConnector[40] = fifoOut[42][2];
              muxOutConnector[41] = fifoOut[43][2];
              muxOutConnector[42] = fifoOut[44][2];
              muxOutConnector[43] = fifoOut[45][2];
              muxOutConnector[44] = fifoOut[46][2];
              muxOutConnector[45] = fifoOut[47][2];
              muxOutConnector[46] = fifoOut[48][2];
              muxOutConnector[47] = fifoOut[49][2];
              muxOutConnector[48] = fifoOut[50][2];
              muxOutConnector[49] = fifoOut[51][2];
              muxOutConnector[50] = fifoOut[26][1];
              muxOutConnector[51] = fifoOut[27][1];
       end
       4: begin
              muxOutConnector[0] = fifoOut[7][11];
              muxOutConnector[1] = fifoOut[8][11];
              muxOutConnector[2] = fifoOut[9][11];
              muxOutConnector[3] = fifoOut[10][11];
              muxOutConnector[4] = fifoOut[11][11];
              muxOutConnector[5] = fifoOut[12][11];
              muxOutConnector[6] = fifoOut[13][11];
              muxOutConnector[7] = fifoOut[14][11];
              muxOutConnector[8] = fifoOut[15][11];
              muxOutConnector[9] = fifoOut[16][11];
              muxOutConnector[10] = fifoOut[17][11];
              muxOutConnector[11] = fifoOut[18][11];
              muxOutConnector[12] = fifoOut[19][11];
              muxOutConnector[13] = fifoOut[20][11];
              muxOutConnector[14] = fifoOut[21][11];
              muxOutConnector[15] = fifoOut[22][11];
              muxOutConnector[16] = fifoOut[23][11];
              muxOutConnector[17] = fifoOut[24][11];
              muxOutConnector[18] = fifoOut[25][11];
              muxOutConnector[19] = fifoOut[0][10];
              muxOutConnector[20] = fifoOut[1][10];
              muxOutConnector[21] = fifoOut[2][10];
              muxOutConnector[22] = fifoOut[3][10];
              muxOutConnector[23] = fifoOut[4][10];
              muxOutConnector[24] = fifoOut[5][10];
              muxOutConnector[25] = fifoOut[6][10];
              muxOutConnector[26] = fifoOut[28][2];
              muxOutConnector[27] = fifoOut[29][2];
              muxOutConnector[28] = fifoOut[30][2];
              muxOutConnector[29] = fifoOut[31][2];
              muxOutConnector[30] = fifoOut[32][2];
              muxOutConnector[31] = fifoOut[33][2];
              muxOutConnector[32] = fifoOut[34][2];
              muxOutConnector[33] = fifoOut[35][2];
              muxOutConnector[34] = fifoOut[36][2];
              muxOutConnector[35] = fifoOut[37][2];
              muxOutConnector[36] = fifoOut[38][2];
              muxOutConnector[37] = fifoOut[39][2];
              muxOutConnector[38] = fifoOut[40][2];
              muxOutConnector[39] = fifoOut[41][2];
              muxOutConnector[40] = fifoOut[42][2];
              muxOutConnector[41] = fifoOut[43][2];
              muxOutConnector[42] = fifoOut[44][2];
              muxOutConnector[43] = fifoOut[45][2];
              muxOutConnector[44] = fifoOut[46][2];
              muxOutConnector[45] = fifoOut[47][2];
              muxOutConnector[46] = fifoOut[48][2];
              muxOutConnector[47] = fifoOut[49][2];
              muxOutConnector[48] = fifoOut[50][2];
              muxOutConnector[49] = fifoOut[51][2];
              muxOutConnector[50] = fifoOut[26][1];
              muxOutConnector[51] = fifoOut[27][1];
       end
       5: begin
              muxOutConnector[0] = fifoOut[7][11];
              muxOutConnector[1] = fifoOut[8][11];
              muxOutConnector[2] = fifoOut[9][11];
              muxOutConnector[3] = fifoOut[10][11];
              muxOutConnector[4] = fifoOut[11][11];
              muxOutConnector[5] = fifoOut[12][11];
              muxOutConnector[6] = fifoOut[13][11];
              muxOutConnector[7] = fifoOut[14][11];
              muxOutConnector[8] = fifoOut[15][11];
              muxOutConnector[9] = fifoOut[16][11];
              muxOutConnector[10] = fifoOut[17][11];
              muxOutConnector[11] = fifoOut[18][11];
              muxOutConnector[12] = fifoOut[19][11];
              muxOutConnector[13] = fifoOut[20][11];
              muxOutConnector[14] = fifoOut[21][11];
              muxOutConnector[15] = fifoOut[22][11];
              muxOutConnector[16] = fifoOut[23][11];
              muxOutConnector[17] = fifoOut[24][11];
              muxOutConnector[18] = fifoOut[25][11];
              muxOutConnector[19] = fifoOut[0][10];
              muxOutConnector[20] = fifoOut[1][10];
              muxOutConnector[21] = fifoOut[2][10];
              muxOutConnector[22] = fifoOut[3][10];
              muxOutConnector[23] = fifoOut[4][10];
              muxOutConnector[24] = fifoOut[5][10];
              muxOutConnector[25] = fifoOut[6][10];
              muxOutConnector[26] = fifoOut[28][2];
              muxOutConnector[27] = fifoOut[29][2];
              muxOutConnector[28] = fifoOut[30][2];
              muxOutConnector[29] = fifoOut[31][2];
              muxOutConnector[30] = fifoOut[32][2];
              muxOutConnector[31] = fifoOut[33][2];
              muxOutConnector[32] = fifoOut[34][2];
              muxOutConnector[33] = fifoOut[35][2];
              muxOutConnector[34] = fifoOut[36][2];
              muxOutConnector[35] = fifoOut[37][2];
              muxOutConnector[36] = fifoOut[38][2];
              muxOutConnector[37] = fifoOut[39][2];
              muxOutConnector[38] = fifoOut[40][2];
              muxOutConnector[39] = fifoOut[41][2];
              muxOutConnector[40] = fifoOut[42][2];
              muxOutConnector[41] = fifoOut[43][2];
              muxOutConnector[42] = fifoOut[44][2];
              muxOutConnector[43] = fifoOut[45][2];
              muxOutConnector[44] = fifoOut[46][2];
              muxOutConnector[45] = fifoOut[47][2];
              muxOutConnector[46] = fifoOut[48][2];
              muxOutConnector[47] = fifoOut[49][2];
              muxOutConnector[48] = fifoOut[50][2];
              muxOutConnector[49] = fifoOut[51][2];
              muxOutConnector[50] = fifoOut[26][1];
              muxOutConnector[51] = fifoOut[27][1];
       end
       6: begin
              muxOutConnector[0] = fifoOut[7][11];
              muxOutConnector[1] = fifoOut[8][11];
              muxOutConnector[2] = fifoOut[9][11];
              muxOutConnector[3] = fifoOut[10][11];
              muxOutConnector[4] = fifoOut[11][11];
              muxOutConnector[5] = fifoOut[12][11];
              muxOutConnector[6] = fifoOut[13][11];
              muxOutConnector[7] = fifoOut[14][11];
              muxOutConnector[8] = fifoOut[15][11];
              muxOutConnector[9] = fifoOut[16][11];
              muxOutConnector[10] = fifoOut[17][11];
              muxOutConnector[11] = fifoOut[18][11];
              muxOutConnector[12] = fifoOut[19][11];
              muxOutConnector[13] = fifoOut[20][11];
              muxOutConnector[14] = fifoOut[21][11];
              muxOutConnector[15] = fifoOut[22][11];
              muxOutConnector[16] = fifoOut[23][11];
              muxOutConnector[17] = fifoOut[24][11];
              muxOutConnector[18] = fifoOut[25][11];
              muxOutConnector[19] = fifoOut[0][10];
              muxOutConnector[20] = fifoOut[1][10];
              muxOutConnector[21] = fifoOut[2][10];
              muxOutConnector[22] = fifoOut[3][10];
              muxOutConnector[23] = fifoOut[4][10];
              muxOutConnector[24] = fifoOut[5][10];
              muxOutConnector[25] = fifoOut[6][10];
              muxOutConnector[26] = fifoOut[28][2];
              muxOutConnector[27] = fifoOut[29][2];
              muxOutConnector[28] = fifoOut[30][2];
              muxOutConnector[29] = fifoOut[31][2];
              muxOutConnector[30] = fifoOut[32][2];
              muxOutConnector[31] = fifoOut[33][2];
              muxOutConnector[32] = fifoOut[34][2];
              muxOutConnector[33] = fifoOut[35][2];
              muxOutConnector[34] = fifoOut[36][2];
              muxOutConnector[35] = fifoOut[37][2];
              muxOutConnector[36] = fifoOut[38][2];
              muxOutConnector[37] = fifoOut[39][2];
              muxOutConnector[38] = fifoOut[40][2];
              muxOutConnector[39] = fifoOut[41][2];
              muxOutConnector[40] = fifoOut[42][2];
              muxOutConnector[41] = fifoOut[43][2];
              muxOutConnector[42] = fifoOut[44][2];
              muxOutConnector[43] = fifoOut[45][2];
              muxOutConnector[44] = fifoOut[46][2];
              muxOutConnector[45] = fifoOut[47][2];
              muxOutConnector[46] = fifoOut[48][2];
              muxOutConnector[47] = fifoOut[49][2];
              muxOutConnector[48] = fifoOut[50][2];
              muxOutConnector[49] = fifoOut[51][2];
              muxOutConnector[50] = fifoOut[26][1];
              muxOutConnector[51] = fifoOut[27][1];
       end
       7: begin
              muxOutConnector[0] = fifoOut[7][11];
              muxOutConnector[1] = fifoOut[8][11];
              muxOutConnector[2] = fifoOut[9][11];
              muxOutConnector[3] = fifoOut[10][11];
              muxOutConnector[4] = fifoOut[11][11];
              muxOutConnector[5] = fifoOut[12][11];
              muxOutConnector[6] = fifoOut[13][11];
              muxOutConnector[7] = fifoOut[14][11];
              muxOutConnector[8] = fifoOut[15][11];
              muxOutConnector[9] = fifoOut[16][11];
              muxOutConnector[10] = fifoOut[17][11];
              muxOutConnector[11] = fifoOut[18][11];
              muxOutConnector[12] = fifoOut[19][11];
              muxOutConnector[13] = fifoOut[20][11];
              muxOutConnector[14] = fifoOut[21][11];
              muxOutConnector[15] = fifoOut[22][11];
              muxOutConnector[16] = fifoOut[23][11];
              muxOutConnector[17] = fifoOut[24][11];
              muxOutConnector[18] = fifoOut[25][11];
              muxOutConnector[19] = fifoOut[0][10];
              muxOutConnector[20] = fifoOut[1][10];
              muxOutConnector[21] = fifoOut[2][10];
              muxOutConnector[22] = fifoOut[3][10];
              muxOutConnector[23] = fifoOut[4][10];
              muxOutConnector[24] = fifoOut[5][10];
              muxOutConnector[25] = fifoOut[6][10];
              muxOutConnector[26] = fifoOut[28][2];
              muxOutConnector[27] = fifoOut[29][2];
              muxOutConnector[28] = fifoOut[30][2];
              muxOutConnector[29] = fifoOut[31][2];
              muxOutConnector[30] = fifoOut[32][2];
              muxOutConnector[31] = fifoOut[33][2];
              muxOutConnector[32] = fifoOut[34][2];
              muxOutConnector[33] = fifoOut[35][2];
              muxOutConnector[34] = fifoOut[36][2];
              muxOutConnector[35] = fifoOut[37][2];
              muxOutConnector[36] = fifoOut[38][2];
              muxOutConnector[37] = fifoOut[39][2];
              muxOutConnector[38] = fifoOut[40][2];
              muxOutConnector[39] = fifoOut[0][6];
              muxOutConnector[40] = fifoOut[1][6];
              muxOutConnector[41] = fifoOut[2][6];
              muxOutConnector[42] = fifoOut[3][6];
              muxOutConnector[43] = fifoOut[4][6];
              muxOutConnector[44] = fifoOut[5][6];
              muxOutConnector[45] = fifoOut[6][6];
              muxOutConnector[46] = fifoOut[7][6];
              muxOutConnector[47] = fifoOut[8][6];
              muxOutConnector[48] = fifoOut[9][6];
              muxOutConnector[49] = fifoOut[10][6];
              muxOutConnector[50] = fifoOut[11][6];
              muxOutConnector[51] = fifoOut[12][6];
       end
       8: begin
              muxOutConnector[0] = fifoOut[7][11];
              muxOutConnector[1] = fifoOut[8][11];
              muxOutConnector[2] = fifoOut[9][11];
              muxOutConnector[3] = fifoOut[10][11];
              muxOutConnector[4] = fifoOut[11][11];
              muxOutConnector[5] = fifoOut[12][11];
              muxOutConnector[6] = fifoOut[13][11];
              muxOutConnector[7] = fifoOut[14][11];
              muxOutConnector[8] = fifoOut[15][11];
              muxOutConnector[9] = fifoOut[16][11];
              muxOutConnector[10] = fifoOut[17][11];
              muxOutConnector[11] = fifoOut[18][11];
              muxOutConnector[12] = fifoOut[19][11];
              muxOutConnector[13] = fifoOut[20][11];
              muxOutConnector[14] = fifoOut[21][11];
              muxOutConnector[15] = fifoOut[22][11];
              muxOutConnector[16] = fifoOut[23][11];
              muxOutConnector[17] = fifoOut[24][11];
              muxOutConnector[18] = fifoOut[25][11];
              muxOutConnector[19] = fifoOut[0][10];
              muxOutConnector[20] = fifoOut[1][10];
              muxOutConnector[21] = fifoOut[2][10];
              muxOutConnector[22] = fifoOut[3][10];
              muxOutConnector[23] = fifoOut[4][10];
              muxOutConnector[24] = fifoOut[5][10];
              muxOutConnector[25] = fifoOut[6][10];
              muxOutConnector[26] = fifoOut[13][7];
              muxOutConnector[27] = fifoOut[14][7];
              muxOutConnector[28] = fifoOut[15][7];
              muxOutConnector[29] = fifoOut[16][7];
              muxOutConnector[30] = fifoOut[17][7];
              muxOutConnector[31] = fifoOut[18][7];
              muxOutConnector[32] = fifoOut[19][7];
              muxOutConnector[33] = fifoOut[20][7];
              muxOutConnector[34] = fifoOut[21][7];
              muxOutConnector[35] = fifoOut[22][7];
              muxOutConnector[36] = fifoOut[23][7];
              muxOutConnector[37] = fifoOut[24][7];
              muxOutConnector[38] = fifoOut[25][7];
              muxOutConnector[39] = fifoOut[0][6];
              muxOutConnector[40] = fifoOut[1][6];
              muxOutConnector[41] = fifoOut[2][6];
              muxOutConnector[42] = fifoOut[3][6];
              muxOutConnector[43] = fifoOut[4][6];
              muxOutConnector[44] = fifoOut[5][6];
              muxOutConnector[45] = fifoOut[6][6];
              muxOutConnector[46] = fifoOut[7][6];
              muxOutConnector[47] = fifoOut[8][6];
              muxOutConnector[48] = fifoOut[9][6];
              muxOutConnector[49] = fifoOut[10][6];
              muxOutConnector[50] = fifoOut[11][6];
              muxOutConnector[51] = fifoOut[12][6];
       end
       9: begin
              muxOutConnector[0] = fifoOut[7][11];
              muxOutConnector[1] = fifoOut[8][11];
              muxOutConnector[2] = fifoOut[9][11];
              muxOutConnector[3] = fifoOut[10][11];
              muxOutConnector[4] = fifoOut[11][11];
              muxOutConnector[5] = fifoOut[12][11];
              muxOutConnector[6] = fifoOut[13][11];
              muxOutConnector[7] = fifoOut[14][11];
              muxOutConnector[8] = fifoOut[15][11];
              muxOutConnector[9] = fifoOut[16][11];
              muxOutConnector[10] = fifoOut[17][11];
              muxOutConnector[11] = fifoOut[18][11];
              muxOutConnector[12] = fifoOut[19][11];
              muxOutConnector[13] = fifoOut[20][11];
              muxOutConnector[14] = fifoOut[21][11];
              muxOutConnector[15] = fifoOut[22][11];
              muxOutConnector[16] = fifoOut[23][11];
              muxOutConnector[17] = fifoOut[24][11];
              muxOutConnector[18] = fifoOut[25][11];
              muxOutConnector[19] = fifoOut[0][10];
              muxOutConnector[20] = fifoOut[1][10];
              muxOutConnector[21] = fifoOut[2][10];
              muxOutConnector[22] = fifoOut[3][10];
              muxOutConnector[23] = fifoOut[4][10];
              muxOutConnector[24] = fifoOut[5][10];
              muxOutConnector[25] = fifoOut[6][10];
              muxOutConnector[26] = fifoOut[13][7];
              muxOutConnector[27] = fifoOut[14][7];
              muxOutConnector[28] = fifoOut[15][7];
              muxOutConnector[29] = fifoOut[16][7];
              muxOutConnector[30] = fifoOut[17][7];
              muxOutConnector[31] = fifoOut[18][7];
              muxOutConnector[32] = fifoOut[19][7];
              muxOutConnector[33] = fifoOut[20][7];
              muxOutConnector[34] = fifoOut[21][7];
              muxOutConnector[35] = fifoOut[22][7];
              muxOutConnector[36] = fifoOut[23][7];
              muxOutConnector[37] = fifoOut[24][7];
              muxOutConnector[38] = fifoOut[25][7];
              muxOutConnector[39] = fifoOut[0][6];
              muxOutConnector[40] = fifoOut[1][6];
              muxOutConnector[41] = fifoOut[2][6];
              muxOutConnector[42] = fifoOut[3][6];
              muxOutConnector[43] = fifoOut[4][6];
              muxOutConnector[44] = fifoOut[5][6];
              muxOutConnector[45] = fifoOut[6][6];
              muxOutConnector[46] = fifoOut[7][6];
              muxOutConnector[47] = fifoOut[8][6];
              muxOutConnector[48] = fifoOut[9][6];
              muxOutConnector[49] = fifoOut[10][6];
              muxOutConnector[50] = fifoOut[11][6];
              muxOutConnector[51] = fifoOut[12][6];
       end
       10: begin
              muxOutConnector[0] = fifoOut[7][11];
              muxOutConnector[1] = fifoOut[8][11];
              muxOutConnector[2] = fifoOut[9][11];
              muxOutConnector[3] = fifoOut[10][11];
              muxOutConnector[4] = fifoOut[11][11];
              muxOutConnector[5] = fifoOut[12][11];
              muxOutConnector[6] = fifoOut[13][11];
              muxOutConnector[7] = fifoOut[14][11];
              muxOutConnector[8] = fifoOut[15][11];
              muxOutConnector[9] = fifoOut[16][11];
              muxOutConnector[10] = fifoOut[17][11];
              muxOutConnector[11] = fifoOut[18][11];
              muxOutConnector[12] = fifoOut[19][11];
              muxOutConnector[13] = fifoOut[20][11];
              muxOutConnector[14] = fifoOut[21][11];
              muxOutConnector[15] = fifoOut[22][11];
              muxOutConnector[16] = fifoOut[23][11];
              muxOutConnector[17] = fifoOut[24][11];
              muxOutConnector[18] = fifoOut[25][11];
              muxOutConnector[19] = fifoOut[0][10];
              muxOutConnector[20] = fifoOut[1][10];
              muxOutConnector[21] = fifoOut[2][10];
              muxOutConnector[22] = fifoOut[3][10];
              muxOutConnector[23] = fifoOut[4][10];
              muxOutConnector[24] = fifoOut[5][10];
              muxOutConnector[25] = fifoOut[6][10];
              muxOutConnector[26] = fifoOut[13][7];
              muxOutConnector[27] = fifoOut[14][7];
              muxOutConnector[28] = fifoOut[15][7];
              muxOutConnector[29] = fifoOut[16][7];
              muxOutConnector[30] = fifoOut[17][7];
              muxOutConnector[31] = fifoOut[18][7];
              muxOutConnector[32] = fifoOut[19][7];
              muxOutConnector[33] = fifoOut[20][7];
              muxOutConnector[34] = fifoOut[21][7];
              muxOutConnector[35] = fifoOut[22][7];
              muxOutConnector[36] = fifoOut[23][7];
              muxOutConnector[37] = fifoOut[24][7];
              muxOutConnector[38] = fifoOut[25][7];
              muxOutConnector[39] = fifoOut[0][6];
              muxOutConnector[40] = fifoOut[1][6];
              muxOutConnector[41] = fifoOut[2][6];
              muxOutConnector[42] = fifoOut[3][6];
              muxOutConnector[43] = fifoOut[4][6];
              muxOutConnector[44] = fifoOut[5][6];
              muxOutConnector[45] = fifoOut[6][6];
              muxOutConnector[46] = fifoOut[7][6];
              muxOutConnector[47] = fifoOut[8][6];
              muxOutConnector[48] = fifoOut[9][6];
              muxOutConnector[49] = fifoOut[10][6];
              muxOutConnector[50] = fifoOut[11][6];
              muxOutConnector[51] = fifoOut[12][6];
       end
       11: begin
              muxOutConnector[0] = fifoOut[7][11];
              muxOutConnector[1] = fifoOut[8][11];
              muxOutConnector[2] = fifoOut[9][11];
              muxOutConnector[3] = fifoOut[10][11];
              muxOutConnector[4] = fifoOut[11][11];
              muxOutConnector[5] = fifoOut[12][11];
              muxOutConnector[6] = fifoOut[13][11];
              muxOutConnector[7] = fifoOut[14][11];
              muxOutConnector[8] = fifoOut[15][11];
              muxOutConnector[9] = fifoOut[16][11];
              muxOutConnector[10] = fifoOut[41][10];
              muxOutConnector[11] = fifoOut[42][10];
              muxOutConnector[12] = fifoOut[43][10];
              muxOutConnector[13] = fifoOut[44][10];
              muxOutConnector[14] = fifoOut[45][10];
              muxOutConnector[15] = fifoOut[46][10];
              muxOutConnector[16] = fifoOut[47][10];
              muxOutConnector[17] = fifoOut[48][10];
              muxOutConnector[18] = fifoOut[49][10];
              muxOutConnector[19] = fifoOut[50][10];
              muxOutConnector[20] = fifoOut[51][10];
              muxOutConnector[21] = fifoOut[26][9];
              muxOutConnector[22] = fifoOut[27][9];
              muxOutConnector[23] = fifoOut[28][9];
              muxOutConnector[24] = fifoOut[29][9];
              muxOutConnector[25] = fifoOut[30][9];
              muxOutConnector[26] = fifoOut[13][7];
              muxOutConnector[27] = fifoOut[14][7];
              muxOutConnector[28] = fifoOut[15][7];
              muxOutConnector[29] = fifoOut[16][7];
              muxOutConnector[30] = fifoOut[17][7];
              muxOutConnector[31] = fifoOut[18][7];
              muxOutConnector[32] = fifoOut[19][7];
              muxOutConnector[33] = fifoOut[20][7];
              muxOutConnector[34] = fifoOut[21][7];
              muxOutConnector[35] = fifoOut[22][7];
              muxOutConnector[36] = fifoOut[23][7];
              muxOutConnector[37] = fifoOut[24][7];
              muxOutConnector[38] = fifoOut[25][7];
              muxOutConnector[39] = fifoOut[0][6];
              muxOutConnector[40] = fifoOut[1][6];
              muxOutConnector[41] = fifoOut[2][6];
              muxOutConnector[42] = fifoOut[3][6];
              muxOutConnector[43] = fifoOut[4][6];
              muxOutConnector[44] = fifoOut[5][6];
              muxOutConnector[45] = fifoOut[6][6];
              muxOutConnector[46] = fifoOut[7][6];
              muxOutConnector[47] = fifoOut[8][6];
              muxOutConnector[48] = fifoOut[9][6];
              muxOutConnector[49] = fifoOut[10][6];
              muxOutConnector[50] = fifoOut[11][6];
              muxOutConnector[51] = fifoOut[12][6];
       end
       12: begin
              muxOutConnector[0] = fifoOut[31][10];
              muxOutConnector[1] = fifoOut[32][10];
              muxOutConnector[2] = fifoOut[33][10];
              muxOutConnector[3] = fifoOut[34][10];
              muxOutConnector[4] = fifoOut[35][10];
              muxOutConnector[5] = fifoOut[36][10];
              muxOutConnector[6] = fifoOut[37][10];
              muxOutConnector[7] = fifoOut[38][10];
              muxOutConnector[8] = fifoOut[39][10];
              muxOutConnector[9] = fifoOut[40][10];
              muxOutConnector[10] = fifoOut[41][10];
              muxOutConnector[11] = fifoOut[42][10];
              muxOutConnector[12] = fifoOut[43][10];
              muxOutConnector[13] = fifoOut[44][10];
              muxOutConnector[14] = fifoOut[45][10];
              muxOutConnector[15] = fifoOut[46][10];
              muxOutConnector[16] = fifoOut[47][10];
              muxOutConnector[17] = fifoOut[48][10];
              muxOutConnector[18] = fifoOut[49][10];
              muxOutConnector[19] = fifoOut[50][10];
              muxOutConnector[20] = fifoOut[51][10];
              muxOutConnector[21] = fifoOut[26][9];
              muxOutConnector[22] = fifoOut[27][9];
              muxOutConnector[23] = fifoOut[28][9];
              muxOutConnector[24] = fifoOut[29][9];
              muxOutConnector[25] = fifoOut[30][9];
              muxOutConnector[26] = fifoOut[13][7];
              muxOutConnector[27] = fifoOut[14][7];
              muxOutConnector[28] = fifoOut[15][7];
              muxOutConnector[29] = fifoOut[16][7];
              muxOutConnector[30] = fifoOut[17][7];
              muxOutConnector[31] = fifoOut[18][7];
              muxOutConnector[32] = fifoOut[19][7];
              muxOutConnector[33] = fifoOut[20][7];
              muxOutConnector[34] = fifoOut[21][7];
              muxOutConnector[35] = fifoOut[22][7];
              muxOutConnector[36] = fifoOut[23][7];
              muxOutConnector[37] = fifoOut[24][7];
              muxOutConnector[38] = fifoOut[25][7];
              muxOutConnector[39] = fifoOut[0][6];
              muxOutConnector[40] = fifoOut[1][6];
              muxOutConnector[41] = fifoOut[2][6];
              muxOutConnector[42] = fifoOut[3][6];
              muxOutConnector[43] = fifoOut[4][6];
              muxOutConnector[44] = fifoOut[5][6];
              muxOutConnector[45] = fifoOut[6][6];
              muxOutConnector[46] = fifoOut[7][6];
              muxOutConnector[47] = fifoOut[8][6];
              muxOutConnector[48] = fifoOut[9][6];
              muxOutConnector[49] = fifoOut[10][6];
              muxOutConnector[50] = fifoOut[11][6];
              muxOutConnector[51] = fifoOut[12][6];
       end
       13: begin
              muxOutConnector[0] = fifoOut[31][10];
              muxOutConnector[1] = fifoOut[32][10];
              muxOutConnector[2] = fifoOut[33][10];
              muxOutConnector[3] = fifoOut[34][10];
              muxOutConnector[4] = fifoOut[35][10];
              muxOutConnector[5] = fifoOut[36][10];
              muxOutConnector[6] = fifoOut[37][10];
              muxOutConnector[7] = fifoOut[38][10];
              muxOutConnector[8] = fifoOut[39][10];
              muxOutConnector[9] = fifoOut[40][10];
              muxOutConnector[10] = fifoOut[41][10];
              muxOutConnector[11] = fifoOut[42][10];
              muxOutConnector[12] = fifoOut[43][10];
              muxOutConnector[13] = fifoOut[44][10];
              muxOutConnector[14] = fifoOut[45][10];
              muxOutConnector[15] = fifoOut[46][10];
              muxOutConnector[16] = fifoOut[47][10];
              muxOutConnector[17] = fifoOut[48][10];
              muxOutConnector[18] = fifoOut[49][10];
              muxOutConnector[19] = fifoOut[50][10];
              muxOutConnector[20] = fifoOut[51][10];
              muxOutConnector[21] = fifoOut[26][9];
              muxOutConnector[22] = fifoOut[27][9];
              muxOutConnector[23] = fifoOut[28][9];
              muxOutConnector[24] = fifoOut[29][9];
              muxOutConnector[25] = fifoOut[30][9];
              muxOutConnector[26] = fifoOut[13][7];
              muxOutConnector[27] = fifoOut[14][7];
              muxOutConnector[28] = fifoOut[15][7];
              muxOutConnector[29] = fifoOut[16][7];
              muxOutConnector[30] = fifoOut[17][7];
              muxOutConnector[31] = fifoOut[18][7];
              muxOutConnector[32] = fifoOut[19][7];
              muxOutConnector[33] = fifoOut[20][7];
              muxOutConnector[34] = fifoOut[21][7];
              muxOutConnector[35] = fifoOut[22][7];
              muxOutConnector[36] = fifoOut[23][7];
              muxOutConnector[37] = fifoOut[24][7];
              muxOutConnector[38] = fifoOut[25][7];
              muxOutConnector[39] = fifoOut[0][6];
              muxOutConnector[40] = fifoOut[1][6];
              muxOutConnector[41] = fifoOut[2][6];
              muxOutConnector[42] = fifoOut[3][6];
              muxOutConnector[43] = fifoOut[4][6];
              muxOutConnector[44] = fifoOut[5][6];
              muxOutConnector[45] = fifoOut[6][6];
              muxOutConnector[46] = fifoOut[7][6];
              muxOutConnector[47] = fifoOut[8][6];
              muxOutConnector[48] = fifoOut[9][6];
              muxOutConnector[49] = fifoOut[10][6];
              muxOutConnector[50] = fifoOut[11][6];
              muxOutConnector[51] = fifoOut[12][6];
       end
       14: begin
              muxOutConnector[0] = fifoOut[31][10];
              muxOutConnector[1] = fifoOut[32][10];
              muxOutConnector[2] = fifoOut[33][10];
              muxOutConnector[3] = fifoOut[34][10];
              muxOutConnector[4] = fifoOut[35][10];
              muxOutConnector[5] = fifoOut[36][10];
              muxOutConnector[6] = fifoOut[37][10];
              muxOutConnector[7] = fifoOut[38][10];
              muxOutConnector[8] = fifoOut[39][10];
              muxOutConnector[9] = fifoOut[40][10];
              muxOutConnector[10] = fifoOut[41][10];
              muxOutConnector[11] = fifoOut[42][10];
              muxOutConnector[12] = fifoOut[43][10];
              muxOutConnector[13] = fifoOut[44][10];
              muxOutConnector[14] = fifoOut[45][10];
              muxOutConnector[15] = fifoOut[46][10];
              muxOutConnector[16] = fifoOut[47][10];
              muxOutConnector[17] = fifoOut[48][10];
              muxOutConnector[18] = fifoOut[49][10];
              muxOutConnector[19] = fifoOut[50][10];
              muxOutConnector[20] = fifoOut[51][10];
              muxOutConnector[21] = fifoOut[26][9];
              muxOutConnector[22] = fifoOut[27][9];
              muxOutConnector[23] = fifoOut[28][9];
              muxOutConnector[24] = fifoOut[29][9];
              muxOutConnector[25] = fifoOut[30][9];
              muxOutConnector[26] = fifoOut[13][7];
              muxOutConnector[27] = fifoOut[14][7];
              muxOutConnector[28] = fifoOut[15][7];
              muxOutConnector[29] = fifoOut[16][7];
              muxOutConnector[30] = fifoOut[17][7];
              muxOutConnector[31] = fifoOut[18][7];
              muxOutConnector[32] = fifoOut[19][7];
              muxOutConnector[33] = fifoOut[20][7];
              muxOutConnector[34] = fifoOut[21][7];
              muxOutConnector[35] = fifoOut[22][7];
              muxOutConnector[36] = fifoOut[23][7];
              muxOutConnector[37] = fifoOut[24][7];
              muxOutConnector[38] = fifoOut[25][7];
              muxOutConnector[39] = fifoOut[0][6];
              muxOutConnector[40] = fifoOut[1][6];
              muxOutConnector[41] = fifoOut[2][6];
              muxOutConnector[42] = fifoOut[3][6];
              muxOutConnector[43] = fifoOut[4][6];
              muxOutConnector[44] = fifoOut[5][6];
              muxOutConnector[45] = fifoOut[6][6];
              muxOutConnector[46] = fifoOut[7][6];
              muxOutConnector[47] = fifoOut[8][6];
              muxOutConnector[48] = fifoOut[9][6];
              muxOutConnector[49] = fifoOut[10][6];
              muxOutConnector[50] = fifoOut[11][6];
              muxOutConnector[51] = fifoOut[12][6];
       end
       15: begin
              muxOutConnector[0] = fifoOut[31][10];
              muxOutConnector[1] = fifoOut[32][10];
              muxOutConnector[2] = fifoOut[33][10];
              muxOutConnector[3] = fifoOut[34][10];
              muxOutConnector[4] = fifoOut[35][10];
              muxOutConnector[5] = fifoOut[36][10];
              muxOutConnector[6] = fifoOut[37][10];
              muxOutConnector[7] = fifoOut[38][10];
              muxOutConnector[8] = fifoOut[39][10];
              muxOutConnector[9] = fifoOut[40][10];
              muxOutConnector[10] = fifoOut[0][14];
              muxOutConnector[11] = fifoOut[1][14];
              muxOutConnector[12] = fifoOut[2][14];
              muxOutConnector[13] = fifoOut[3][14];
              muxOutConnector[14] = fifoOut[4][14];
              muxOutConnector[15] = fifoOut[5][14];
              muxOutConnector[16] = fifoOut[6][14];
              muxOutConnector[17] = fifoOut[7][14];
              muxOutConnector[18] = fifoOut[8][14];
              muxOutConnector[19] = fifoOut[9][14];
              muxOutConnector[20] = fifoOut[10][14];
              muxOutConnector[21] = fifoOut[11][14];
              muxOutConnector[22] = fifoOut[12][14];
              muxOutConnector[23] = fifoOut[13][14];
              muxOutConnector[24] = fifoOut[14][14];
              muxOutConnector[25] = fifoOut[15][14];
              muxOutConnector[26] = fifoOut[13][7];
              muxOutConnector[27] = fifoOut[14][7];
              muxOutConnector[28] = fifoOut[15][7];
              muxOutConnector[29] = fifoOut[16][7];
              muxOutConnector[30] = fifoOut[17][7];
              muxOutConnector[31] = fifoOut[18][7];
              muxOutConnector[32] = fifoOut[19][7];
              muxOutConnector[33] = fifoOut[20][7];
              muxOutConnector[34] = fifoOut[21][7];
              muxOutConnector[35] = fifoOut[22][7];
              muxOutConnector[36] = fifoOut[23][7];
              muxOutConnector[37] = fifoOut[24][7];
              muxOutConnector[38] = fifoOut[25][7];
              muxOutConnector[39] = fifoOut[0][6];
              muxOutConnector[40] = fifoOut[1][6];
              muxOutConnector[41] = fifoOut[2][6];
              muxOutConnector[42] = fifoOut[3][6];
              muxOutConnector[43] = fifoOut[4][6];
              muxOutConnector[44] = fifoOut[5][6];
              muxOutConnector[45] = fifoOut[6][6];
              muxOutConnector[46] = fifoOut[7][6];
              muxOutConnector[47] = fifoOut[8][6];
              muxOutConnector[48] = fifoOut[9][6];
              muxOutConnector[49] = fifoOut[10][6];
              muxOutConnector[50] = fifoOut[11][6];
              muxOutConnector[51] = fifoOut[12][6];
       end
       16: begin
              muxOutConnector[0] = fifoOut[16][15];
              muxOutConnector[1] = fifoOut[17][15];
              muxOutConnector[2] = fifoOut[18][15];
              muxOutConnector[3] = fifoOut[19][15];
              muxOutConnector[4] = fifoOut[20][15];
              muxOutConnector[5] = fifoOut[21][15];
              muxOutConnector[6] = fifoOut[22][15];
              muxOutConnector[7] = fifoOut[23][15];
              muxOutConnector[8] = fifoOut[24][15];
              muxOutConnector[9] = fifoOut[25][15];
              muxOutConnector[10] = fifoOut[0][14];
              muxOutConnector[11] = fifoOut[1][14];
              muxOutConnector[12] = fifoOut[2][14];
              muxOutConnector[13] = fifoOut[3][14];
              muxOutConnector[14] = fifoOut[4][14];
              muxOutConnector[15] = fifoOut[5][14];
              muxOutConnector[16] = fifoOut[6][14];
              muxOutConnector[17] = fifoOut[7][14];
              muxOutConnector[18] = fifoOut[8][14];
              muxOutConnector[19] = fifoOut[9][14];
              muxOutConnector[20] = fifoOut[10][14];
              muxOutConnector[21] = fifoOut[11][14];
              muxOutConnector[22] = fifoOut[12][14];
              muxOutConnector[23] = fifoOut[13][14];
              muxOutConnector[24] = fifoOut[14][14];
              muxOutConnector[25] = fifoOut[15][14];
              muxOutConnector[26] = fifoOut[13][7];
              muxOutConnector[27] = fifoOut[14][7];
              muxOutConnector[28] = fifoOut[15][7];
              muxOutConnector[29] = fifoOut[16][7];
              muxOutConnector[30] = fifoOut[17][7];
              muxOutConnector[31] = fifoOut[18][7];
              muxOutConnector[32] = fifoOut[19][7];
              muxOutConnector[33] = fifoOut[20][7];
              muxOutConnector[34] = fifoOut[21][7];
              muxOutConnector[35] = fifoOut[22][7];
              muxOutConnector[36] = fifoOut[23][7];
              muxOutConnector[37] = fifoOut[24][7];
              muxOutConnector[38] = fifoOut[25][7];
              muxOutConnector[39] = fifoOut[0][6];
              muxOutConnector[40] = fifoOut[1][6];
              muxOutConnector[41] = fifoOut[2][6];
              muxOutConnector[42] = fifoOut[3][6];
              muxOutConnector[43] = fifoOut[4][6];
              muxOutConnector[44] = fifoOut[5][6];
              muxOutConnector[45] = fifoOut[6][6];
              muxOutConnector[46] = fifoOut[7][6];
              muxOutConnector[47] = fifoOut[8][6];
              muxOutConnector[48] = fifoOut[9][6];
              muxOutConnector[49] = fifoOut[10][6];
              muxOutConnector[50] = fifoOut[11][6];
              muxOutConnector[51] = fifoOut[12][6];
       end
       17: begin
              muxOutConnector[0] = fifoOut[16][15];
              muxOutConnector[1] = fifoOut[17][15];
              muxOutConnector[2] = fifoOut[18][15];
              muxOutConnector[3] = fifoOut[19][15];
              muxOutConnector[4] = fifoOut[20][15];
              muxOutConnector[5] = fifoOut[21][15];
              muxOutConnector[6] = fifoOut[22][15];
              muxOutConnector[7] = fifoOut[23][15];
              muxOutConnector[8] = fifoOut[24][15];
              muxOutConnector[9] = fifoOut[25][15];
              muxOutConnector[10] = fifoOut[0][14];
              muxOutConnector[11] = fifoOut[1][14];
              muxOutConnector[12] = fifoOut[2][14];
              muxOutConnector[13] = fifoOut[3][14];
              muxOutConnector[14] = fifoOut[4][14];
              muxOutConnector[15] = fifoOut[5][14];
              muxOutConnector[16] = fifoOut[6][14];
              muxOutConnector[17] = fifoOut[7][14];
              muxOutConnector[18] = fifoOut[8][14];
              muxOutConnector[19] = fifoOut[9][14];
              muxOutConnector[20] = fifoOut[10][14];
              muxOutConnector[21] = fifoOut[11][14];
              muxOutConnector[22] = fifoOut[12][14];
              muxOutConnector[23] = fifoOut[13][14];
              muxOutConnector[24] = fifoOut[14][14];
              muxOutConnector[25] = fifoOut[15][14];
              muxOutConnector[26] = fifoOut[13][7];
              muxOutConnector[27] = fifoOut[14][7];
              muxOutConnector[28] = fifoOut[15][7];
              muxOutConnector[29] = fifoOut[16][7];
              muxOutConnector[30] = fifoOut[17][7];
              muxOutConnector[31] = fifoOut[18][7];
              muxOutConnector[32] = fifoOut[19][7];
              muxOutConnector[33] = fifoOut[20][7];
              muxOutConnector[34] = fifoOut[21][7];
              muxOutConnector[35] = fifoOut[22][7];
              muxOutConnector[36] = fifoOut[23][7];
              muxOutConnector[37] = fifoOut[24][7];
              muxOutConnector[38] = fifoOut[25][7];
              muxOutConnector[39] = fifoOut[0][6];
              muxOutConnector[40] = fifoOut[1][6];
              muxOutConnector[41] = fifoOut[2][6];
              muxOutConnector[42] = fifoOut[3][6];
              muxOutConnector[43] = fifoOut[4][6];
              muxOutConnector[44] = fifoOut[5][6];
              muxOutConnector[45] = fifoOut[6][6];
              muxOutConnector[46] = fifoOut[7][6];
              muxOutConnector[47] = fifoOut[8][6];
              muxOutConnector[48] = fifoOut[9][6];
              muxOutConnector[49] = fifoOut[10][6];
              muxOutConnector[50] = fifoOut[11][6];
              muxOutConnector[51] = fifoOut[12][6];
       end
       18: begin
              muxOutConnector[0] = fifoOut[16][15];
              muxOutConnector[1] = fifoOut[17][15];
              muxOutConnector[2] = fifoOut[18][15];
              muxOutConnector[3] = fifoOut[19][15];
              muxOutConnector[4] = fifoOut[20][15];
              muxOutConnector[5] = fifoOut[21][15];
              muxOutConnector[6] = fifoOut[22][15];
              muxOutConnector[7] = fifoOut[23][15];
              muxOutConnector[8] = fifoOut[24][15];
              muxOutConnector[9] = fifoOut[25][15];
              muxOutConnector[10] = fifoOut[0][14];
              muxOutConnector[11] = fifoOut[1][14];
              muxOutConnector[12] = fifoOut[2][14];
              muxOutConnector[13] = fifoOut[3][14];
              muxOutConnector[14] = fifoOut[4][14];
              muxOutConnector[15] = fifoOut[5][14];
              muxOutConnector[16] = fifoOut[6][14];
              muxOutConnector[17] = fifoOut[7][14];
              muxOutConnector[18] = fifoOut[8][14];
              muxOutConnector[19] = fifoOut[9][14];
              muxOutConnector[20] = fifoOut[10][14];
              muxOutConnector[21] = fifoOut[11][14];
              muxOutConnector[22] = fifoOut[12][14];
              muxOutConnector[23] = fifoOut[13][14];
              muxOutConnector[24] = fifoOut[14][14];
              muxOutConnector[25] = fifoOut[15][14];
              muxOutConnector[26] = fifoOut[13][7];
              muxOutConnector[27] = fifoOut[14][7];
              muxOutConnector[28] = fifoOut[15][7];
              muxOutConnector[29] = fifoOut[16][7];
              muxOutConnector[30] = fifoOut[17][7];
              muxOutConnector[31] = fifoOut[18][7];
              muxOutConnector[32] = fifoOut[19][7];
              muxOutConnector[33] = fifoOut[20][7];
              muxOutConnector[34] = fifoOut[21][7];
              muxOutConnector[35] = fifoOut[22][7];
              muxOutConnector[36] = fifoOut[23][7];
              muxOutConnector[37] = fifoOut[24][7];
              muxOutConnector[38] = fifoOut[25][7];
              muxOutConnector[39] = fifoOut[0][6];
              muxOutConnector[40] = fifoOut[1][6];
              muxOutConnector[41] = fifoOut[2][6];
              muxOutConnector[42] = fifoOut[3][6];
              muxOutConnector[43] = fifoOut[4][6];
              muxOutConnector[44] = fifoOut[5][6];
              muxOutConnector[45] = fifoOut[6][6];
              muxOutConnector[46] = fifoOut[7][6];
              muxOutConnector[47] = fifoOut[8][6];
              muxOutConnector[48] = fifoOut[9][6];
              muxOutConnector[49] = fifoOut[10][6];
              muxOutConnector[50] = fifoOut[11][6];
              muxOutConnector[51] = fifoOut[12][6];
       end
       19: begin
              muxOutConnector[0] = fifoOut[16][15];
              muxOutConnector[1] = fifoOut[17][15];
              muxOutConnector[2] = fifoOut[18][15];
              muxOutConnector[3] = fifoOut[19][15];
              muxOutConnector[4] = fifoOut[20][15];
              muxOutConnector[5] = fifoOut[21][15];
              muxOutConnector[6] = fifoOut[22][15];
              muxOutConnector[7] = fifoOut[23][15];
              muxOutConnector[8] = fifoOut[24][15];
              muxOutConnector[9] = fifoOut[25][15];
              muxOutConnector[10] = fifoOut[0][14];
              muxOutConnector[11] = fifoOut[1][14];
              muxOutConnector[12] = fifoOut[2][14];
              muxOutConnector[13] = fifoOut[3][14];
              muxOutConnector[14] = fifoOut[4][14];
              muxOutConnector[15] = fifoOut[5][14];
              muxOutConnector[16] = fifoOut[6][14];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[13][7];
              muxOutConnector[27] = fifoOut[14][7];
              muxOutConnector[28] = fifoOut[15][7];
              muxOutConnector[29] = fifoOut[16][7];
              muxOutConnector[30] = fifoOut[17][7];
              muxOutConnector[31] = fifoOut[18][7];
              muxOutConnector[32] = fifoOut[19][7];
              muxOutConnector[33] = fifoOut[20][7];
              muxOutConnector[34] = fifoOut[21][7];
              muxOutConnector[35] = fifoOut[22][7];
              muxOutConnector[36] = fifoOut[23][7];
              muxOutConnector[37] = fifoOut[24][7];
              muxOutConnector[38] = fifoOut[25][7];
              muxOutConnector[39] = fifoOut[0][6];
              muxOutConnector[40] = fifoOut[1][6];
              muxOutConnector[41] = fifoOut[2][6];
              muxOutConnector[42] = fifoOut[3][6];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
