`timescale 1ns / 1ps
module LMem1To0_511_circ6_combined_ys_yu_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        rxIn,
        load_input_en,
        iteration_0_indicator,
        feedback_en,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter r_lower = 32;
parameter c = 17;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input load_input_en;
input iteration_0_indicator;
input [ADDRESSWIDTH-1:0]unloadAddress;
input feedback_en;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input [ r_lower * w - 1 : 0 ] rxIn; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
wire [w-1:0]rxInConnector[r_lower-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

generate
    for (k=0;k<r_lower;k=k+1)begin:assign_rx
        assign rxInConnector[k] = rxIn[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            if(feedback_en)begin
                 fifoOut[i][0] <= fifoOut[i][c-1];
            end
            else if(load_input_en)begin
                 if(i < r_lower)begin
                   fifoOut[i][0] = rxInConnector[i];
                 end
                 else begin
                   fifoOut[i][0] = maxVal;
                 end
            end
            else begin
                 fifoOut[i][0] <= ly0InConnector[i];
            end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
       0: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = fifoOut[21][2][w-1];
              unloadMuxOut[27] = fifoOut[22][2][w-1];
              unloadMuxOut[28] = fifoOut[23][2][w-1];
              unloadMuxOut[29] = fifoOut[24][2][w-1];
              unloadMuxOut[30] = fifoOut[25][2][w-1];
              unloadMuxOut[31] = fifoOut[0][1][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[1][2][w-1];
              unloadMuxOut[1] = fifoOut[2][2][w-1];
              unloadMuxOut[2] = fifoOut[3][2][w-1];
              unloadMuxOut[3] = fifoOut[4][2][w-1];
              unloadMuxOut[4] = fifoOut[5][2][w-1];
              unloadMuxOut[5] = fifoOut[6][2][w-1];
              unloadMuxOut[6] = fifoOut[7][2][w-1];
              unloadMuxOut[7] = fifoOut[8][2][w-1];
              unloadMuxOut[8] = fifoOut[9][2][w-1];
              unloadMuxOut[9] = fifoOut[10][2][w-1];
              unloadMuxOut[10] = fifoOut[11][2][w-1];
              unloadMuxOut[11] = fifoOut[12][2][w-1];
              unloadMuxOut[12] = fifoOut[13][2][w-1];
              unloadMuxOut[13] = fifoOut[14][2][w-1];
              unloadMuxOut[14] = fifoOut[15][2][w-1];
              unloadMuxOut[15] = fifoOut[16][2][w-1];
              unloadMuxOut[16] = fifoOut[17][2][w-1];
              unloadMuxOut[17] = fifoOut[18][2][w-1];
              unloadMuxOut[18] = fifoOut[19][2][w-1];
              unloadMuxOut[19] = fifoOut[20][2][w-1];
              unloadMuxOut[20] = fifoOut[21][2][w-1];
              unloadMuxOut[21] = fifoOut[22][2][w-1];
              unloadMuxOut[22] = fifoOut[23][2][w-1];
              unloadMuxOut[23] = fifoOut[24][2][w-1];
              unloadMuxOut[24] = fifoOut[25][2][w-1];
              unloadMuxOut[25] = fifoOut[0][1][w-1];
              unloadMuxOut[26] = fifoOut[1][1][w-1];
              unloadMuxOut[27] = fifoOut[2][1][w-1];
              unloadMuxOut[28] = fifoOut[3][1][w-1];
              unloadMuxOut[29] = fifoOut[4][1][w-1];
              unloadMuxOut[30] = fifoOut[5][1][w-1];
              unloadMuxOut[31] = fifoOut[6][1][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[7][2][w-1];
              unloadMuxOut[1] = fifoOut[8][2][w-1];
              unloadMuxOut[2] = fifoOut[9][2][w-1];
              unloadMuxOut[3] = fifoOut[26][15][w-1];
              unloadMuxOut[4] = fifoOut[27][15][w-1];
              unloadMuxOut[5] = fifoOut[28][15][w-1];
              unloadMuxOut[6] = fifoOut[29][15][w-1];
              unloadMuxOut[7] = fifoOut[30][15][w-1];
              unloadMuxOut[8] = fifoOut[31][15][w-1];
              unloadMuxOut[9] = fifoOut[32][15][w-1];
              unloadMuxOut[10] = fifoOut[33][15][w-1];
              unloadMuxOut[11] = fifoOut[34][15][w-1];
              unloadMuxOut[12] = fifoOut[35][15][w-1];
              unloadMuxOut[13] = fifoOut[36][15][w-1];
              unloadMuxOut[14] = fifoOut[37][15][w-1];
              unloadMuxOut[15] = fifoOut[38][15][w-1];
              unloadMuxOut[16] = fifoOut[39][15][w-1];
              unloadMuxOut[17] = fifoOut[40][15][w-1];
              unloadMuxOut[18] = fifoOut[41][15][w-1];
              unloadMuxOut[19] = fifoOut[42][15][w-1];
              unloadMuxOut[20] = fifoOut[43][15][w-1];
              unloadMuxOut[21] = fifoOut[44][15][w-1];
              unloadMuxOut[22] = fifoOut[45][15][w-1];
              unloadMuxOut[23] = fifoOut[46][15][w-1];
              unloadMuxOut[24] = fifoOut[47][15][w-1];
              unloadMuxOut[25] = fifoOut[48][15][w-1];
              unloadMuxOut[26] = fifoOut[49][15][w-1];
              unloadMuxOut[27] = fifoOut[50][15][w-1];
              unloadMuxOut[28] = fifoOut[51][15][w-1];
              unloadMuxOut[29] = fifoOut[26][14][w-1];
              unloadMuxOut[30] = fifoOut[27][14][w-1];
              unloadMuxOut[31] = fifoOut[28][14][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[29][15][w-1];
              unloadMuxOut[1] = fifoOut[30][15][w-1];
              unloadMuxOut[2] = fifoOut[31][15][w-1];
              unloadMuxOut[3] = fifoOut[32][15][w-1];
              unloadMuxOut[4] = fifoOut[33][15][w-1];
              unloadMuxOut[5] = fifoOut[34][15][w-1];
              unloadMuxOut[6] = fifoOut[35][15][w-1];
              unloadMuxOut[7] = fifoOut[36][15][w-1];
              unloadMuxOut[8] = fifoOut[37][15][w-1];
              unloadMuxOut[9] = fifoOut[38][15][w-1];
              unloadMuxOut[10] = fifoOut[39][15][w-1];
              unloadMuxOut[11] = fifoOut[40][15][w-1];
              unloadMuxOut[12] = fifoOut[41][15][w-1];
              unloadMuxOut[13] = fifoOut[42][15][w-1];
              unloadMuxOut[14] = fifoOut[43][15][w-1];
              unloadMuxOut[15] = fifoOut[44][15][w-1];
              unloadMuxOut[16] = fifoOut[45][15][w-1];
              unloadMuxOut[17] = fifoOut[46][15][w-1];
              unloadMuxOut[18] = fifoOut[47][15][w-1];
              unloadMuxOut[19] = fifoOut[48][15][w-1];
              unloadMuxOut[20] = fifoOut[49][15][w-1];
              unloadMuxOut[21] = fifoOut[50][15][w-1];
              unloadMuxOut[22] = fifoOut[51][15][w-1];
              unloadMuxOut[23] = fifoOut[26][14][w-1];
              unloadMuxOut[24] = fifoOut[27][14][w-1];
              unloadMuxOut[25] = fifoOut[28][14][w-1];
              unloadMuxOut[26] = fifoOut[29][14][w-1];
              unloadMuxOut[27] = fifoOut[30][14][w-1];
              unloadMuxOut[28] = fifoOut[31][14][w-1];
              unloadMuxOut[29] = fifoOut[32][14][w-1];
              unloadMuxOut[30] = fifoOut[33][14][w-1];
              unloadMuxOut[31] = fifoOut[34][14][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[35][15][w-1];
              unloadMuxOut[1] = fifoOut[36][15][w-1];
              unloadMuxOut[2] = fifoOut[37][15][w-1];
              unloadMuxOut[3] = fifoOut[38][15][w-1];
              unloadMuxOut[4] = fifoOut[39][15][w-1];
              unloadMuxOut[5] = fifoOut[40][15][w-1];
              unloadMuxOut[6] = fifoOut[41][15][w-1];
              unloadMuxOut[7] = fifoOut[42][15][w-1];
              unloadMuxOut[8] = fifoOut[43][15][w-1];
              unloadMuxOut[9] = fifoOut[44][15][w-1];
              unloadMuxOut[10] = fifoOut[45][15][w-1];
              unloadMuxOut[11] = fifoOut[46][15][w-1];
              unloadMuxOut[12] = fifoOut[47][15][w-1];
              unloadMuxOut[13] = fifoOut[48][15][w-1];
              unloadMuxOut[14] = fifoOut[49][15][w-1];
              unloadMuxOut[15] = fifoOut[50][15][w-1];
              unloadMuxOut[16] = fifoOut[51][15][w-1];
              unloadMuxOut[17] = fifoOut[26][14][w-1];
              unloadMuxOut[18] = fifoOut[27][14][w-1];
              unloadMuxOut[19] = fifoOut[28][14][w-1];
              unloadMuxOut[20] = fifoOut[29][14][w-1];
              unloadMuxOut[21] = fifoOut[30][14][w-1];
              unloadMuxOut[22] = fifoOut[31][14][w-1];
              unloadMuxOut[23] = fifoOut[32][14][w-1];
              unloadMuxOut[24] = fifoOut[33][14][w-1];
              unloadMuxOut[25] = fifoOut[34][14][w-1];
              unloadMuxOut[26] = fifoOut[35][14][w-1];
              unloadMuxOut[27] = fifoOut[36][14][w-1];
              unloadMuxOut[28] = fifoOut[37][14][w-1];
              unloadMuxOut[29] = fifoOut[38][14][w-1];
              unloadMuxOut[30] = fifoOut[39][14][w-1];
              unloadMuxOut[31] = fifoOut[40][14][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[41][15][w-1];
              unloadMuxOut[1] = fifoOut[42][15][w-1];
              unloadMuxOut[2] = fifoOut[43][15][w-1];
              unloadMuxOut[3] = fifoOut[44][15][w-1];
              unloadMuxOut[4] = fifoOut[45][15][w-1];
              unloadMuxOut[5] = fifoOut[46][15][w-1];
              unloadMuxOut[6] = fifoOut[47][15][w-1];
              unloadMuxOut[7] = fifoOut[48][15][w-1];
              unloadMuxOut[8] = fifoOut[49][15][w-1];
              unloadMuxOut[9] = fifoOut[50][15][w-1];
              unloadMuxOut[10] = fifoOut[51][15][w-1];
              unloadMuxOut[11] = fifoOut[26][14][w-1];
              unloadMuxOut[12] = fifoOut[27][14][w-1];
              unloadMuxOut[13] = fifoOut[28][14][w-1];
              unloadMuxOut[14] = fifoOut[29][14][w-1];
              unloadMuxOut[15] = fifoOut[30][14][w-1];
              unloadMuxOut[16] = fifoOut[31][14][w-1];
              unloadMuxOut[17] = fifoOut[32][14][w-1];
              unloadMuxOut[18] = fifoOut[33][14][w-1];
              unloadMuxOut[19] = fifoOut[34][14][w-1];
              unloadMuxOut[20] = fifoOut[35][14][w-1];
              unloadMuxOut[21] = fifoOut[36][14][w-1];
              unloadMuxOut[22] = fifoOut[37][14][w-1];
              unloadMuxOut[23] = fifoOut[38][14][w-1];
              unloadMuxOut[24] = fifoOut[39][14][w-1];
              unloadMuxOut[25] = fifoOut[40][14][w-1];
              unloadMuxOut[26] = fifoOut[41][14][w-1];
              unloadMuxOut[27] = fifoOut[42][14][w-1];
              unloadMuxOut[28] = fifoOut[43][14][w-1];
              unloadMuxOut[29] = fifoOut[44][14][w-1];
              unloadMuxOut[30] = fifoOut[45][14][w-1];
              unloadMuxOut[31] = fifoOut[46][14][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[47][15][w-1];
              unloadMuxOut[1] = fifoOut[48][15][w-1];
              unloadMuxOut[2] = fifoOut[49][15][w-1];
              unloadMuxOut[3] = fifoOut[50][15][w-1];
              unloadMuxOut[4] = fifoOut[51][15][w-1];
              unloadMuxOut[5] = fifoOut[26][14][w-1];
              unloadMuxOut[6] = fifoOut[27][14][w-1];
              unloadMuxOut[7] = fifoOut[28][14][w-1];
              unloadMuxOut[8] = fifoOut[29][14][w-1];
              unloadMuxOut[9] = fifoOut[30][14][w-1];
              unloadMuxOut[10] = fifoOut[31][14][w-1];
              unloadMuxOut[11] = fifoOut[32][14][w-1];
              unloadMuxOut[12] = fifoOut[33][14][w-1];
              unloadMuxOut[13] = fifoOut[34][14][w-1];
              unloadMuxOut[14] = fifoOut[35][14][w-1];
              unloadMuxOut[15] = fifoOut[36][14][w-1];
              unloadMuxOut[16] = fifoOut[37][14][w-1];
              unloadMuxOut[17] = fifoOut[38][14][w-1];
              unloadMuxOut[18] = fifoOut[39][14][w-1];
              unloadMuxOut[19] = fifoOut[40][14][w-1];
              unloadMuxOut[20] = fifoOut[41][14][w-1];
              unloadMuxOut[21] = fifoOut[42][14][w-1];
              unloadMuxOut[22] = fifoOut[43][14][w-1];
              unloadMuxOut[23] = fifoOut[44][14][w-1];
              unloadMuxOut[24] = fifoOut[45][14][w-1];
              unloadMuxOut[25] = fifoOut[46][14][w-1];
              unloadMuxOut[26] = fifoOut[47][14][w-1];
              unloadMuxOut[27] = fifoOut[48][14][w-1];
              unloadMuxOut[28] = fifoOut[49][14][w-1];
              unloadMuxOut[29] = fifoOut[50][14][w-1];
              unloadMuxOut[30] = fifoOut[51][14][w-1];
              unloadMuxOut[31] = fifoOut[26][13][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[27][14][w-1];
              unloadMuxOut[1] = fifoOut[28][14][w-1];
              unloadMuxOut[2] = fifoOut[29][14][w-1];
              unloadMuxOut[3] = fifoOut[30][14][w-1];
              unloadMuxOut[4] = fifoOut[31][14][w-1];
              unloadMuxOut[5] = fifoOut[32][14][w-1];
              unloadMuxOut[6] = fifoOut[33][14][w-1];
              unloadMuxOut[7] = fifoOut[34][14][w-1];
              unloadMuxOut[8] = fifoOut[35][14][w-1];
              unloadMuxOut[9] = fifoOut[36][14][w-1];
              unloadMuxOut[10] = fifoOut[37][14][w-1];
              unloadMuxOut[11] = fifoOut[38][14][w-1];
              unloadMuxOut[12] = fifoOut[39][14][w-1];
              unloadMuxOut[13] = fifoOut[40][14][w-1];
              unloadMuxOut[14] = fifoOut[41][14][w-1];
              unloadMuxOut[15] = fifoOut[42][14][w-1];
              unloadMuxOut[16] = fifoOut[43][14][w-1];
              unloadMuxOut[17] = fifoOut[44][14][w-1];
              unloadMuxOut[18] = fifoOut[45][14][w-1];
              unloadMuxOut[19] = fifoOut[46][14][w-1];
              unloadMuxOut[20] = fifoOut[47][14][w-1];
              unloadMuxOut[21] = fifoOut[48][14][w-1];
              unloadMuxOut[22] = fifoOut[49][14][w-1];
              unloadMuxOut[23] = fifoOut[50][14][w-1];
              unloadMuxOut[24] = fifoOut[51][14][w-1];
              unloadMuxOut[25] = fifoOut[26][13][w-1];
              unloadMuxOut[26] = fifoOut[27][13][w-1];
              unloadMuxOut[27] = fifoOut[28][13][w-1];
              unloadMuxOut[28] = fifoOut[29][13][w-1];
              unloadMuxOut[29] = fifoOut[30][13][w-1];
              unloadMuxOut[30] = fifoOut[31][13][w-1];
              unloadMuxOut[31] = fifoOut[32][13][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[33][14][w-1];
              unloadMuxOut[1] = fifoOut[34][14][w-1];
              unloadMuxOut[2] = fifoOut[35][14][w-1];
              unloadMuxOut[3] = fifoOut[36][14][w-1];
              unloadMuxOut[4] = fifoOut[37][14][w-1];
              unloadMuxOut[5] = fifoOut[38][14][w-1];
              unloadMuxOut[6] = fifoOut[39][14][w-1];
              unloadMuxOut[7] = fifoOut[40][14][w-1];
              unloadMuxOut[8] = fifoOut[41][14][w-1];
              unloadMuxOut[9] = fifoOut[42][14][w-1];
              unloadMuxOut[10] = fifoOut[43][14][w-1];
              unloadMuxOut[11] = fifoOut[44][14][w-1];
              unloadMuxOut[12] = fifoOut[45][14][w-1];
              unloadMuxOut[13] = fifoOut[46][14][w-1];
              unloadMuxOut[14] = fifoOut[47][14][w-1];
              unloadMuxOut[15] = fifoOut[48][14][w-1];
              unloadMuxOut[16] = fifoOut[49][14][w-1];
              unloadMuxOut[17] = fifoOut[50][14][w-1];
              unloadMuxOut[18] = fifoOut[51][14][w-1];
              unloadMuxOut[19] = fifoOut[26][13][w-1];
              unloadMuxOut[20] = fifoOut[27][13][w-1];
              unloadMuxOut[21] = fifoOut[28][13][w-1];
              unloadMuxOut[22] = fifoOut[29][13][w-1];
              unloadMuxOut[23] = fifoOut[30][13][w-1];
              unloadMuxOut[24] = fifoOut[31][13][w-1];
              unloadMuxOut[25] = fifoOut[32][13][w-1];
              unloadMuxOut[26] = fifoOut[33][13][w-1];
              unloadMuxOut[27] = fifoOut[34][13][w-1];
              unloadMuxOut[28] = fifoOut[35][13][w-1];
              unloadMuxOut[29] = fifoOut[36][13][w-1];
              unloadMuxOut[30] = fifoOut[37][13][w-1];
              unloadMuxOut[31] = fifoOut[38][13][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[39][14][w-1];
              unloadMuxOut[1] = fifoOut[40][14][w-1];
              unloadMuxOut[2] = fifoOut[41][14][w-1];
              unloadMuxOut[3] = fifoOut[42][14][w-1];
              unloadMuxOut[4] = fifoOut[43][14][w-1];
              unloadMuxOut[5] = fifoOut[44][14][w-1];
              unloadMuxOut[6] = fifoOut[45][14][w-1];
              unloadMuxOut[7] = fifoOut[46][14][w-1];
              unloadMuxOut[8] = fifoOut[47][14][w-1];
              unloadMuxOut[9] = fifoOut[48][14][w-1];
              unloadMuxOut[10] = fifoOut[49][14][w-1];
              unloadMuxOut[11] = fifoOut[50][14][w-1];
              unloadMuxOut[12] = fifoOut[51][14][w-1];
              unloadMuxOut[13] = fifoOut[26][13][w-1];
              unloadMuxOut[14] = fifoOut[27][13][w-1];
              unloadMuxOut[15] = fifoOut[28][13][w-1];
              unloadMuxOut[16] = fifoOut[29][13][w-1];
              unloadMuxOut[17] = fifoOut[30][13][w-1];
              unloadMuxOut[18] = fifoOut[31][13][w-1];
              unloadMuxOut[19] = fifoOut[32][13][w-1];
              unloadMuxOut[20] = fifoOut[33][13][w-1];
              unloadMuxOut[21] = fifoOut[34][13][w-1];
              unloadMuxOut[22] = fifoOut[35][13][w-1];
              unloadMuxOut[23] = fifoOut[36][13][w-1];
              unloadMuxOut[24] = fifoOut[37][13][w-1];
              unloadMuxOut[25] = fifoOut[38][13][w-1];
              unloadMuxOut[26] = fifoOut[39][13][w-1];
              unloadMuxOut[27] = fifoOut[40][13][w-1];
              unloadMuxOut[28] = fifoOut[41][13][w-1];
              unloadMuxOut[29] = fifoOut[42][13][w-1];
              unloadMuxOut[30] = fifoOut[43][13][w-1];
              unloadMuxOut[31] = fifoOut[44][13][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[45][14][w-1];
              unloadMuxOut[1] = fifoOut[46][14][w-1];
              unloadMuxOut[2] = fifoOut[47][14][w-1];
              unloadMuxOut[3] = fifoOut[48][14][w-1];
              unloadMuxOut[4] = fifoOut[49][14][w-1];
              unloadMuxOut[5] = fifoOut[50][14][w-1];
              unloadMuxOut[6] = fifoOut[51][14][w-1];
              unloadMuxOut[7] = fifoOut[26][13][w-1];
              unloadMuxOut[8] = fifoOut[27][13][w-1];
              unloadMuxOut[9] = fifoOut[28][13][w-1];
              unloadMuxOut[10] = fifoOut[29][13][w-1];
              unloadMuxOut[11] = fifoOut[30][13][w-1];
              unloadMuxOut[12] = fifoOut[31][13][w-1];
              unloadMuxOut[13] = fifoOut[32][13][w-1];
              unloadMuxOut[14] = fifoOut[33][13][w-1];
              unloadMuxOut[15] = fifoOut[34][13][w-1];
              unloadMuxOut[16] = fifoOut[35][13][w-1];
              unloadMuxOut[17] = fifoOut[36][13][w-1];
              unloadMuxOut[18] = fifoOut[37][13][w-1];
              unloadMuxOut[19] = fifoOut[38][13][w-1];
              unloadMuxOut[20] = fifoOut[39][13][w-1];
              unloadMuxOut[21] = fifoOut[40][13][w-1];
              unloadMuxOut[22] = fifoOut[41][13][w-1];
              unloadMuxOut[23] = fifoOut[42][13][w-1];
              unloadMuxOut[24] = fifoOut[43][13][w-1];
              unloadMuxOut[25] = fifoOut[44][13][w-1];
              unloadMuxOut[26] = fifoOut[45][13][w-1];
              unloadMuxOut[27] = fifoOut[46][13][w-1];
              unloadMuxOut[28] = fifoOut[47][13][w-1];
              unloadMuxOut[29] = fifoOut[48][13][w-1];
              unloadMuxOut[30] = fifoOut[49][13][w-1];
              unloadMuxOut[31] = fifoOut[50][13][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[51][14][w-1];
              unloadMuxOut[1] = fifoOut[26][13][w-1];
              unloadMuxOut[2] = fifoOut[27][13][w-1];
              unloadMuxOut[3] = fifoOut[28][13][w-1];
              unloadMuxOut[4] = fifoOut[29][13][w-1];
              unloadMuxOut[5] = fifoOut[30][13][w-1];
              unloadMuxOut[6] = fifoOut[31][13][w-1];
              unloadMuxOut[7] = fifoOut[32][13][w-1];
              unloadMuxOut[8] = fifoOut[33][13][w-1];
              unloadMuxOut[9] = fifoOut[34][13][w-1];
              unloadMuxOut[10] = fifoOut[35][13][w-1];
              unloadMuxOut[11] = fifoOut[36][13][w-1];
              unloadMuxOut[12] = fifoOut[37][13][w-1];
              unloadMuxOut[13] = fifoOut[38][13][w-1];
              unloadMuxOut[14] = fifoOut[39][13][w-1];
              unloadMuxOut[15] = fifoOut[40][13][w-1];
              unloadMuxOut[16] = fifoOut[41][13][w-1];
              unloadMuxOut[17] = fifoOut[42][13][w-1];
              unloadMuxOut[18] = fifoOut[43][13][w-1];
              unloadMuxOut[19] = fifoOut[44][13][w-1];
              unloadMuxOut[20] = fifoOut[45][13][w-1];
              unloadMuxOut[21] = fifoOut[46][13][w-1];
              unloadMuxOut[22] = fifoOut[47][13][w-1];
              unloadMuxOut[23] = fifoOut[48][13][w-1];
              unloadMuxOut[24] = fifoOut[49][13][w-1];
              unloadMuxOut[25] = fifoOut[50][13][w-1];
              unloadMuxOut[26] = fifoOut[51][13][w-1];
              unloadMuxOut[27] = fifoOut[26][12][w-1];
              unloadMuxOut[28] = fifoOut[27][12][w-1];
              unloadMuxOut[29] = fifoOut[28][12][w-1];
              unloadMuxOut[30] = fifoOut[29][12][w-1];
              unloadMuxOut[31] = fifoOut[30][12][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[31][13][w-1];
              unloadMuxOut[1] = fifoOut[32][13][w-1];
              unloadMuxOut[2] = fifoOut[33][13][w-1];
              unloadMuxOut[3] = fifoOut[34][13][w-1];
              unloadMuxOut[4] = fifoOut[35][13][w-1];
              unloadMuxOut[5] = fifoOut[36][13][w-1];
              unloadMuxOut[6] = fifoOut[37][13][w-1];
              unloadMuxOut[7] = fifoOut[38][13][w-1];
              unloadMuxOut[8] = fifoOut[39][13][w-1];
              unloadMuxOut[9] = fifoOut[40][13][w-1];
              unloadMuxOut[10] = fifoOut[41][13][w-1];
              unloadMuxOut[11] = fifoOut[42][13][w-1];
              unloadMuxOut[12] = fifoOut[43][13][w-1];
              unloadMuxOut[13] = fifoOut[44][13][w-1];
              unloadMuxOut[14] = fifoOut[45][13][w-1];
              unloadMuxOut[15] = fifoOut[46][13][w-1];
              unloadMuxOut[16] = fifoOut[47][13][w-1];
              unloadMuxOut[17] = fifoOut[48][13][w-1];
              unloadMuxOut[18] = fifoOut[49][13][w-1];
              unloadMuxOut[19] = fifoOut[50][13][w-1];
              unloadMuxOut[20] = fifoOut[51][13][w-1];
              unloadMuxOut[21] = fifoOut[26][12][w-1];
              unloadMuxOut[22] = fifoOut[27][12][w-1];
              unloadMuxOut[23] = fifoOut[28][12][w-1];
              unloadMuxOut[24] = fifoOut[29][12][w-1];
              unloadMuxOut[25] = fifoOut[30][12][w-1];
              unloadMuxOut[26] = fifoOut[31][12][w-1];
              unloadMuxOut[27] = fifoOut[32][12][w-1];
              unloadMuxOut[28] = fifoOut[33][12][w-1];
              unloadMuxOut[29] = fifoOut[34][12][w-1];
              unloadMuxOut[30] = fifoOut[35][12][w-1];
              unloadMuxOut[31] = fifoOut[36][12][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[37][13][w-1];
              unloadMuxOut[1] = fifoOut[38][13][w-1];
              unloadMuxOut[2] = fifoOut[39][13][w-1];
              unloadMuxOut[3] = fifoOut[40][13][w-1];
              unloadMuxOut[4] = fifoOut[41][13][w-1];
              unloadMuxOut[5] = fifoOut[42][13][w-1];
              unloadMuxOut[6] = fifoOut[10][2][w-1];
              unloadMuxOut[7] = fifoOut[11][2][w-1];
              unloadMuxOut[8] = fifoOut[12][2][w-1];
              unloadMuxOut[9] = fifoOut[13][2][w-1];
              unloadMuxOut[10] = fifoOut[14][2][w-1];
              unloadMuxOut[11] = fifoOut[15][2][w-1];
              unloadMuxOut[12] = fifoOut[16][2][w-1];
              unloadMuxOut[13] = fifoOut[17][2][w-1];
              unloadMuxOut[14] = fifoOut[18][2][w-1];
              unloadMuxOut[15] = fifoOut[19][2][w-1];
              unloadMuxOut[16] = fifoOut[20][2][w-1];
              unloadMuxOut[17] = fifoOut[21][2][w-1];
              unloadMuxOut[18] = fifoOut[22][2][w-1];
              unloadMuxOut[19] = fifoOut[23][2][w-1];
              unloadMuxOut[20] = fifoOut[24][2][w-1];
              unloadMuxOut[21] = fifoOut[25][2][w-1];
              unloadMuxOut[22] = fifoOut[0][1][w-1];
              unloadMuxOut[23] = fifoOut[1][1][w-1];
              unloadMuxOut[24] = fifoOut[2][1][w-1];
              unloadMuxOut[25] = fifoOut[3][1][w-1];
              unloadMuxOut[26] = fifoOut[4][1][w-1];
              unloadMuxOut[27] = fifoOut[5][1][w-1];
              unloadMuxOut[28] = fifoOut[6][1][w-1];
              unloadMuxOut[29] = fifoOut[7][1][w-1];
              unloadMuxOut[30] = fifoOut[8][1][w-1];
              unloadMuxOut[31] = fifoOut[9][1][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[10][2][w-1];
              unloadMuxOut[1] = fifoOut[11][2][w-1];
              unloadMuxOut[2] = fifoOut[12][2][w-1];
              unloadMuxOut[3] = fifoOut[13][2][w-1];
              unloadMuxOut[4] = fifoOut[14][2][w-1];
              unloadMuxOut[5] = fifoOut[15][2][w-1];
              unloadMuxOut[6] = fifoOut[16][2][w-1];
              unloadMuxOut[7] = fifoOut[17][2][w-1];
              unloadMuxOut[8] = fifoOut[18][2][w-1];
              unloadMuxOut[9] = fifoOut[19][2][w-1];
              unloadMuxOut[10] = fifoOut[20][2][w-1];
              unloadMuxOut[11] = fifoOut[21][2][w-1];
              unloadMuxOut[12] = fifoOut[22][2][w-1];
              unloadMuxOut[13] = fifoOut[23][2][w-1];
              unloadMuxOut[14] = fifoOut[24][2][w-1];
              unloadMuxOut[15] = fifoOut[25][2][w-1];
              unloadMuxOut[16] = fifoOut[0][1][w-1];
              unloadMuxOut[17] = fifoOut[1][1][w-1];
              unloadMuxOut[18] = fifoOut[2][1][w-1];
              unloadMuxOut[19] = fifoOut[3][1][w-1];
              unloadMuxOut[20] = fifoOut[4][1][w-1];
              unloadMuxOut[21] = fifoOut[5][1][w-1];
              unloadMuxOut[22] = fifoOut[6][1][w-1];
              unloadMuxOut[23] = fifoOut[7][1][w-1];
              unloadMuxOut[24] = fifoOut[8][1][w-1];
              unloadMuxOut[25] = fifoOut[9][1][w-1];
              unloadMuxOut[26] = fifoOut[10][1][w-1];
              unloadMuxOut[27] = fifoOut[11][1][w-1];
              unloadMuxOut[28] = fifoOut[12][1][w-1];
              unloadMuxOut[29] = fifoOut[13][1][w-1];
              unloadMuxOut[30] = fifoOut[14][1][w-1];
              unloadMuxOut[31] = fifoOut[15][1][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[16][2][w-1];
              unloadMuxOut[1] = fifoOut[17][2][w-1];
              unloadMuxOut[2] = fifoOut[18][2][w-1];
              unloadMuxOut[3] = fifoOut[19][2][w-1];
              unloadMuxOut[4] = fifoOut[20][2][w-1];
              unloadMuxOut[5] = fifoOut[21][2][w-1];
              unloadMuxOut[6] = fifoOut[22][2][w-1];
              unloadMuxOut[7] = fifoOut[23][2][w-1];
              unloadMuxOut[8] = fifoOut[24][2][w-1];
              unloadMuxOut[9] = fifoOut[25][2][w-1];
              unloadMuxOut[10] = fifoOut[0][1][w-1];
              unloadMuxOut[11] = fifoOut[1][1][w-1];
              unloadMuxOut[12] = fifoOut[2][1][w-1];
              unloadMuxOut[13] = fifoOut[3][1][w-1];
              unloadMuxOut[14] = fifoOut[4][1][w-1];
              unloadMuxOut[15] = fifoOut[5][1][w-1];
              unloadMuxOut[16] = fifoOut[6][1][w-1];
              unloadMuxOut[17] = fifoOut[7][1][w-1];
              unloadMuxOut[18] = fifoOut[8][1][w-1];
              unloadMuxOut[19] = fifoOut[9][1][w-1];
              unloadMuxOut[20] = fifoOut[10][1][w-1];
              unloadMuxOut[21] = fifoOut[11][1][w-1];
              unloadMuxOut[22] = fifoOut[12][1][w-1];
              unloadMuxOut[23] = fifoOut[13][1][w-1];
              unloadMuxOut[24] = fifoOut[14][1][w-1];
              unloadMuxOut[25] = fifoOut[15][1][w-1];
              unloadMuxOut[26] = fifoOut[16][1][w-1];
              unloadMuxOut[27] = fifoOut[17][1][w-1];
              unloadMuxOut[28] = fifoOut[18][1][w-1];
              unloadMuxOut[29] = fifoOut[19][1][w-1];
              unloadMuxOut[30] = fifoOut[20][1][w-1];
              unloadMuxOut[31] = fifoOut[21][1][w-1];
       end
       16: begin
              unloadMuxOut[0] = fifoOut[22][2][w-1];
              unloadMuxOut[1] = fifoOut[23][2][w-1];
              unloadMuxOut[2] = fifoOut[24][2][w-1];
              unloadMuxOut[3] = fifoOut[25][2][w-1];
              unloadMuxOut[4] = fifoOut[0][1][w-1];
              unloadMuxOut[5] = fifoOut[1][1][w-1];
              unloadMuxOut[6] = fifoOut[2][1][w-1];
              unloadMuxOut[7] = fifoOut[3][1][w-1];
              unloadMuxOut[8] = fifoOut[4][1][w-1];
              unloadMuxOut[9] = fifoOut[5][1][w-1];
              unloadMuxOut[10] = fifoOut[6][1][w-1];
              unloadMuxOut[11] = fifoOut[7][1][w-1];
              unloadMuxOut[12] = fifoOut[8][1][w-1];
              unloadMuxOut[13] = fifoOut[9][1][w-1];
              unloadMuxOut[14] = fifoOut[10][1][w-1];
              unloadMuxOut[15] = fifoOut[11][1][w-1];
              unloadMuxOut[16] = fifoOut[12][1][w-1];
              unloadMuxOut[17] = fifoOut[13][1][w-1];
              unloadMuxOut[18] = fifoOut[14][1][w-1];
              unloadMuxOut[19] = fifoOut[15][1][w-1];
              unloadMuxOut[20] = fifoOut[16][1][w-1];
              unloadMuxOut[21] = fifoOut[17][1][w-1];
              unloadMuxOut[22] = fifoOut[18][1][w-1];
              unloadMuxOut[23] = fifoOut[19][1][w-1];
              unloadMuxOut[24] = fifoOut[20][1][w-1];
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0; 
             end
       end
    endcase //unload case end
    case(iteration_0_indicator)
       0: begin
         case(rd_address_case)
         0: begin
              muxOutConnector[0] = fifoOut[21][2];
              muxOutConnector[1] = fifoOut[22][2];
              muxOutConnector[2] = fifoOut[23][2];
              muxOutConnector[3] = fifoOut[24][2];
              muxOutConnector[4] = fifoOut[25][2];
              muxOutConnector[5] = fifoOut[0][1];
              muxOutConnector[6] = fifoOut[1][1];
              muxOutConnector[7] = fifoOut[2][1];
              muxOutConnector[8] = fifoOut[3][1];
              muxOutConnector[9] = fifoOut[4][1];
              muxOutConnector[10] = fifoOut[5][1];
              muxOutConnector[11] = fifoOut[6][1];
              muxOutConnector[12] = fifoOut[7][1];
              muxOutConnector[13] = fifoOut[8][1];
              muxOutConnector[14] = fifoOut[9][1];
              muxOutConnector[15] = fifoOut[10][1];
              muxOutConnector[16] = fifoOut[11][1];
              muxOutConnector[17] = fifoOut[12][1];
              muxOutConnector[18] = fifoOut[13][1];
              muxOutConnector[19] = fifoOut[14][1];
              muxOutConnector[20] = fifoOut[15][1];
              muxOutConnector[21] = fifoOut[16][1];
              muxOutConnector[22] = fifoOut[17][1];
              muxOutConnector[23] = fifoOut[18][1];
              muxOutConnector[24] = fifoOut[19][1];
              muxOutConnector[25] = fifoOut[20][1];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
         end
         1: begin
              muxOutConnector[0] = fifoOut[21][2];
              muxOutConnector[1] = fifoOut[22][2];
              muxOutConnector[2] = fifoOut[23][2];
              muxOutConnector[3] = fifoOut[24][2];
              muxOutConnector[4] = fifoOut[25][2];
              muxOutConnector[5] = fifoOut[0][1];
              muxOutConnector[6] = fifoOut[1][1];
              muxOutConnector[7] = fifoOut[2][1];
              muxOutConnector[8] = fifoOut[3][1];
              muxOutConnector[9] = fifoOut[4][1];
              muxOutConnector[10] = fifoOut[5][1];
              muxOutConnector[11] = fifoOut[6][1];
              muxOutConnector[12] = fifoOut[7][1];
              muxOutConnector[13] = fifoOut[8][1];
              muxOutConnector[14] = fifoOut[9][1];
              muxOutConnector[15] = fifoOut[26][14];
              muxOutConnector[16] = fifoOut[27][14];
              muxOutConnector[17] = fifoOut[28][14];
              muxOutConnector[18] = fifoOut[29][14];
              muxOutConnector[19] = fifoOut[30][14];
              muxOutConnector[20] = fifoOut[31][14];
              muxOutConnector[21] = fifoOut[32][14];
              muxOutConnector[22] = fifoOut[33][14];
              muxOutConnector[23] = fifoOut[34][14];
              muxOutConnector[24] = fifoOut[35][14];
              muxOutConnector[25] = fifoOut[36][14];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
         end
         2: begin
              muxOutConnector[0] = fifoOut[37][15];
              muxOutConnector[1] = fifoOut[38][15];
              muxOutConnector[2] = fifoOut[39][15];
              muxOutConnector[3] = fifoOut[40][15];
              muxOutConnector[4] = fifoOut[41][15];
              muxOutConnector[5] = fifoOut[42][15];
              muxOutConnector[6] = fifoOut[43][15];
              muxOutConnector[7] = fifoOut[44][15];
              muxOutConnector[8] = fifoOut[45][15];
              muxOutConnector[9] = fifoOut[46][15];
              muxOutConnector[10] = fifoOut[47][15];
              muxOutConnector[11] = fifoOut[48][15];
              muxOutConnector[12] = fifoOut[49][15];
              muxOutConnector[13] = fifoOut[50][15];
              muxOutConnector[14] = fifoOut[51][15];
              muxOutConnector[15] = fifoOut[26][14];
              muxOutConnector[16] = fifoOut[27][14];
              muxOutConnector[17] = fifoOut[28][14];
              muxOutConnector[18] = fifoOut[29][14];
              muxOutConnector[19] = fifoOut[30][14];
              muxOutConnector[20] = fifoOut[31][14];
              muxOutConnector[21] = fifoOut[32][14];
              muxOutConnector[22] = fifoOut[33][14];
              muxOutConnector[23] = fifoOut[34][14];
              muxOutConnector[24] = fifoOut[35][14];
              muxOutConnector[25] = fifoOut[36][14];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
         end
         3: begin
              muxOutConnector[0] = fifoOut[37][15];
              muxOutConnector[1] = fifoOut[38][15];
              muxOutConnector[2] = fifoOut[39][15];
              muxOutConnector[3] = fifoOut[40][15];
              muxOutConnector[4] = fifoOut[41][15];
              muxOutConnector[5] = fifoOut[42][15];
              muxOutConnector[6] = fifoOut[43][15];
              muxOutConnector[7] = fifoOut[44][15];
              muxOutConnector[8] = fifoOut[45][15];
              muxOutConnector[9] = fifoOut[46][15];
              muxOutConnector[10] = fifoOut[47][15];
              muxOutConnector[11] = fifoOut[48][15];
              muxOutConnector[12] = fifoOut[49][15];
              muxOutConnector[13] = fifoOut[50][15];
              muxOutConnector[14] = fifoOut[51][15];
              muxOutConnector[15] = fifoOut[26][14];
              muxOutConnector[16] = fifoOut[27][14];
              muxOutConnector[17] = fifoOut[28][14];
              muxOutConnector[18] = fifoOut[29][14];
              muxOutConnector[19] = fifoOut[30][14];
              muxOutConnector[20] = fifoOut[31][14];
              muxOutConnector[21] = fifoOut[32][14];
              muxOutConnector[22] = fifoOut[33][14];
              muxOutConnector[23] = fifoOut[34][14];
              muxOutConnector[24] = fifoOut[35][14];
              muxOutConnector[25] = fifoOut[36][14];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
         end
         4: begin
              muxOutConnector[0] = fifoOut[37][15];
              muxOutConnector[1] = fifoOut[38][15];
              muxOutConnector[2] = fifoOut[39][15];
              muxOutConnector[3] = fifoOut[40][15];
              muxOutConnector[4] = fifoOut[41][15];
              muxOutConnector[5] = fifoOut[42][15];
              muxOutConnector[6] = fifoOut[43][15];
              muxOutConnector[7] = fifoOut[44][15];
              muxOutConnector[8] = fifoOut[45][15];
              muxOutConnector[9] = fifoOut[46][15];
              muxOutConnector[10] = fifoOut[47][15];
              muxOutConnector[11] = fifoOut[48][15];
              muxOutConnector[12] = fifoOut[49][15];
              muxOutConnector[13] = fifoOut[50][15];
              muxOutConnector[14] = fifoOut[51][15];
              muxOutConnector[15] = fifoOut[26][14];
              muxOutConnector[16] = fifoOut[27][14];
              muxOutConnector[17] = fifoOut[28][14];
              muxOutConnector[18] = fifoOut[29][14];
              muxOutConnector[19] = fifoOut[30][14];
              muxOutConnector[20] = fifoOut[31][14];
              muxOutConnector[21] = fifoOut[32][14];
              muxOutConnector[22] = fifoOut[33][14];
              muxOutConnector[23] = fifoOut[34][14];
              muxOutConnector[24] = fifoOut[35][14];
              muxOutConnector[25] = fifoOut[36][14];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
         end
         5: begin
              muxOutConnector[0] = fifoOut[37][15];
              muxOutConnector[1] = fifoOut[38][15];
              muxOutConnector[2] = fifoOut[39][15];
              muxOutConnector[3] = fifoOut[40][15];
              muxOutConnector[4] = fifoOut[41][15];
              muxOutConnector[5] = fifoOut[42][15];
              muxOutConnector[6] = fifoOut[43][15];
              muxOutConnector[7] = fifoOut[44][15];
              muxOutConnector[8] = fifoOut[45][15];
              muxOutConnector[9] = fifoOut[46][15];
              muxOutConnector[10] = fifoOut[47][15];
              muxOutConnector[11] = fifoOut[48][15];
              muxOutConnector[12] = fifoOut[49][15];
              muxOutConnector[13] = fifoOut[50][15];
              muxOutConnector[14] = fifoOut[51][15];
              muxOutConnector[15] = fifoOut[26][14];
              muxOutConnector[16] = fifoOut[27][14];
              muxOutConnector[17] = fifoOut[28][14];
              muxOutConnector[18] = fifoOut[29][14];
              muxOutConnector[19] = fifoOut[30][14];
              muxOutConnector[20] = fifoOut[31][14];
              muxOutConnector[21] = fifoOut[32][14];
              muxOutConnector[22] = fifoOut[33][14];
              muxOutConnector[23] = fifoOut[34][14];
              muxOutConnector[24] = fifoOut[35][14];
              muxOutConnector[25] = fifoOut[36][14];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
         end
         6: begin
              muxOutConnector[0] = fifoOut[37][15];
              muxOutConnector[1] = fifoOut[38][15];
              muxOutConnector[2] = fifoOut[39][15];
              muxOutConnector[3] = fifoOut[40][15];
              muxOutConnector[4] = fifoOut[41][15];
              muxOutConnector[5] = fifoOut[42][15];
              muxOutConnector[6] = fifoOut[43][15];
              muxOutConnector[7] = fifoOut[44][15];
              muxOutConnector[8] = fifoOut[45][15];
              muxOutConnector[9] = fifoOut[46][15];
              muxOutConnector[10] = fifoOut[47][15];
              muxOutConnector[11] = fifoOut[48][15];
              muxOutConnector[12] = fifoOut[49][15];
              muxOutConnector[13] = fifoOut[50][15];
              muxOutConnector[14] = fifoOut[51][15];
              muxOutConnector[15] = fifoOut[26][14];
              muxOutConnector[16] = fifoOut[27][14];
              muxOutConnector[17] = fifoOut[28][14];
              muxOutConnector[18] = fifoOut[29][14];
              muxOutConnector[19] = fifoOut[30][14];
              muxOutConnector[20] = fifoOut[31][14];
              muxOutConnector[21] = fifoOut[32][14];
              muxOutConnector[22] = fifoOut[33][14];
              muxOutConnector[23] = fifoOut[34][14];
              muxOutConnector[24] = fifoOut[35][14];
              muxOutConnector[25] = fifoOut[36][14];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
         end
         7: begin
              muxOutConnector[0] = fifoOut[37][15];
              muxOutConnector[1] = fifoOut[38][15];
              muxOutConnector[2] = fifoOut[39][15];
              muxOutConnector[3] = fifoOut[40][15];
              muxOutConnector[4] = fifoOut[41][15];
              muxOutConnector[5] = fifoOut[42][15];
              muxOutConnector[6] = fifoOut[43][15];
              muxOutConnector[7] = fifoOut[44][15];
              muxOutConnector[8] = fifoOut[45][15];
              muxOutConnector[9] = fifoOut[46][15];
              muxOutConnector[10] = fifoOut[47][15];
              muxOutConnector[11] = fifoOut[48][15];
              muxOutConnector[12] = fifoOut[49][15];
              muxOutConnector[13] = fifoOut[50][15];
              muxOutConnector[14] = fifoOut[51][15];
              muxOutConnector[15] = fifoOut[26][14];
              muxOutConnector[16] = fifoOut[27][14];
              muxOutConnector[17] = fifoOut[28][14];
              muxOutConnector[18] = fifoOut[29][14];
              muxOutConnector[19] = fifoOut[30][14];
              muxOutConnector[20] = fifoOut[31][14];
              muxOutConnector[21] = fifoOut[32][14];
              muxOutConnector[22] = fifoOut[33][14];
              muxOutConnector[23] = fifoOut[34][14];
              muxOutConnector[24] = fifoOut[35][14];
              muxOutConnector[25] = fifoOut[36][14];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
         end
         8: begin
              muxOutConnector[0] = fifoOut[37][15];
              muxOutConnector[1] = fifoOut[38][15];
              muxOutConnector[2] = fifoOut[39][15];
              muxOutConnector[3] = fifoOut[40][15];
              muxOutConnector[4] = fifoOut[41][15];
              muxOutConnector[5] = fifoOut[42][15];
              muxOutConnector[6] = fifoOut[43][15];
              muxOutConnector[7] = fifoOut[44][15];
              muxOutConnector[8] = fifoOut[45][15];
              muxOutConnector[9] = fifoOut[46][15];
              muxOutConnector[10] = fifoOut[47][15];
              muxOutConnector[11] = fifoOut[48][15];
              muxOutConnector[12] = fifoOut[49][15];
              muxOutConnector[13] = fifoOut[50][15];
              muxOutConnector[14] = fifoOut[51][15];
              muxOutConnector[15] = fifoOut[26][14];
              muxOutConnector[16] = fifoOut[27][14];
              muxOutConnector[17] = fifoOut[28][14];
              muxOutConnector[18] = fifoOut[29][14];
              muxOutConnector[19] = fifoOut[30][14];
              muxOutConnector[20] = fifoOut[31][14];
              muxOutConnector[21] = fifoOut[32][14];
              muxOutConnector[22] = fifoOut[33][14];
              muxOutConnector[23] = fifoOut[34][14];
              muxOutConnector[24] = fifoOut[35][14];
              muxOutConnector[25] = fifoOut[36][14];
              muxOutConnector[26] = fifoOut[33][4];
              muxOutConnector[27] = fifoOut[34][4];
              muxOutConnector[28] = fifoOut[35][4];
              muxOutConnector[29] = fifoOut[36][4];
              muxOutConnector[30] = fifoOut[37][4];
              muxOutConnector[31] = fifoOut[38][4];
              muxOutConnector[32] = fifoOut[39][4];
              muxOutConnector[33] = fifoOut[40][4];
              muxOutConnector[34] = fifoOut[41][4];
              muxOutConnector[35] = fifoOut[42][4];
              muxOutConnector[36] = fifoOut[43][4];
              muxOutConnector[37] = fifoOut[44][4];
              muxOutConnector[38] = fifoOut[45][4];
              muxOutConnector[39] = fifoOut[46][4];
              muxOutConnector[40] = fifoOut[47][4];
              muxOutConnector[41] = fifoOut[48][4];
              muxOutConnector[42] = fifoOut[49][4];
              muxOutConnector[43] = fifoOut[50][4];
              muxOutConnector[44] = fifoOut[51][4];
              muxOutConnector[45] = fifoOut[26][3];
              muxOutConnector[46] = fifoOut[27][3];
              muxOutConnector[47] = fifoOut[28][3];
              muxOutConnector[48] = fifoOut[29][3];
              muxOutConnector[49] = fifoOut[30][3];
              muxOutConnector[50] = fifoOut[31][3];
              muxOutConnector[51] = fifoOut[32][3];
         end
         9: begin
              muxOutConnector[0] = fifoOut[37][15];
              muxOutConnector[1] = fifoOut[38][15];
              muxOutConnector[2] = fifoOut[39][15];
              muxOutConnector[3] = fifoOut[40][15];
              muxOutConnector[4] = fifoOut[41][15];
              muxOutConnector[5] = fifoOut[42][15];
              muxOutConnector[6] = fifoOut[43][15];
              muxOutConnector[7] = fifoOut[44][15];
              muxOutConnector[8] = fifoOut[45][15];
              muxOutConnector[9] = fifoOut[46][15];
              muxOutConnector[10] = fifoOut[47][15];
              muxOutConnector[11] = fifoOut[48][15];
              muxOutConnector[12] = fifoOut[49][15];
              muxOutConnector[13] = fifoOut[50][15];
              muxOutConnector[14] = fifoOut[51][15];
              muxOutConnector[15] = fifoOut[26][14];
              muxOutConnector[16] = fifoOut[27][14];
              muxOutConnector[17] = fifoOut[28][14];
              muxOutConnector[18] = fifoOut[29][14];
              muxOutConnector[19] = fifoOut[30][14];
              muxOutConnector[20] = fifoOut[31][14];
              muxOutConnector[21] = fifoOut[32][14];
              muxOutConnector[22] = fifoOut[33][14];
              muxOutConnector[23] = fifoOut[34][14];
              muxOutConnector[24] = fifoOut[35][14];
              muxOutConnector[25] = fifoOut[36][14];
              muxOutConnector[26] = fifoOut[33][4];
              muxOutConnector[27] = fifoOut[34][4];
              muxOutConnector[28] = fifoOut[35][4];
              muxOutConnector[29] = fifoOut[36][4];
              muxOutConnector[30] = fifoOut[37][4];
              muxOutConnector[31] = fifoOut[38][4];
              muxOutConnector[32] = fifoOut[39][4];
              muxOutConnector[33] = fifoOut[40][4];
              muxOutConnector[34] = fifoOut[41][4];
              muxOutConnector[35] = fifoOut[42][4];
              muxOutConnector[36] = fifoOut[43][4];
              muxOutConnector[37] = fifoOut[44][4];
              muxOutConnector[38] = fifoOut[45][4];
              muxOutConnector[39] = fifoOut[46][4];
              muxOutConnector[40] = fifoOut[47][4];
              muxOutConnector[41] = fifoOut[48][4];
              muxOutConnector[42] = fifoOut[49][4];
              muxOutConnector[43] = fifoOut[50][4];
              muxOutConnector[44] = fifoOut[51][4];
              muxOutConnector[45] = fifoOut[26][3];
              muxOutConnector[46] = fifoOut[27][3];
              muxOutConnector[47] = fifoOut[28][3];
              muxOutConnector[48] = fifoOut[29][3];
              muxOutConnector[49] = fifoOut[30][3];
              muxOutConnector[50] = fifoOut[31][3];
              muxOutConnector[51] = fifoOut[32][3];
         end
         10: begin
              muxOutConnector[0] = fifoOut[37][15];
              muxOutConnector[1] = fifoOut[38][15];
              muxOutConnector[2] = fifoOut[39][15];
              muxOutConnector[3] = fifoOut[40][15];
              muxOutConnector[4] = fifoOut[41][15];
              muxOutConnector[5] = fifoOut[42][15];
              muxOutConnector[6] = fifoOut[43][15];
              muxOutConnector[7] = fifoOut[44][15];
              muxOutConnector[8] = fifoOut[45][15];
              muxOutConnector[9] = fifoOut[46][15];
              muxOutConnector[10] = fifoOut[47][15];
              muxOutConnector[11] = fifoOut[48][15];
              muxOutConnector[12] = fifoOut[49][15];
              muxOutConnector[13] = fifoOut[50][15];
              muxOutConnector[14] = fifoOut[51][15];
              muxOutConnector[15] = fifoOut[26][14];
              muxOutConnector[16] = fifoOut[27][14];
              muxOutConnector[17] = fifoOut[28][14];
              muxOutConnector[18] = fifoOut[29][14];
              muxOutConnector[19] = fifoOut[30][14];
              muxOutConnector[20] = fifoOut[31][14];
              muxOutConnector[21] = fifoOut[32][14];
              muxOutConnector[22] = fifoOut[33][14];
              muxOutConnector[23] = fifoOut[34][14];
              muxOutConnector[24] = fifoOut[35][14];
              muxOutConnector[25] = fifoOut[36][14];
              muxOutConnector[26] = fifoOut[33][4];
              muxOutConnector[27] = fifoOut[34][4];
              muxOutConnector[28] = fifoOut[35][4];
              muxOutConnector[29] = fifoOut[36][4];
              muxOutConnector[30] = fifoOut[37][4];
              muxOutConnector[31] = fifoOut[38][4];
              muxOutConnector[32] = fifoOut[39][4];
              muxOutConnector[33] = fifoOut[40][4];
              muxOutConnector[34] = fifoOut[41][4];
              muxOutConnector[35] = fifoOut[42][4];
              muxOutConnector[36] = fifoOut[43][4];
              muxOutConnector[37] = fifoOut[44][4];
              muxOutConnector[38] = fifoOut[45][4];
              muxOutConnector[39] = fifoOut[46][4];
              muxOutConnector[40] = fifoOut[47][4];
              muxOutConnector[41] = fifoOut[48][4];
              muxOutConnector[42] = fifoOut[49][4];
              muxOutConnector[43] = fifoOut[50][4];
              muxOutConnector[44] = fifoOut[51][4];
              muxOutConnector[45] = fifoOut[26][3];
              muxOutConnector[46] = fifoOut[27][3];
              muxOutConnector[47] = fifoOut[28][3];
              muxOutConnector[48] = fifoOut[29][3];
              muxOutConnector[49] = fifoOut[30][3];
              muxOutConnector[50] = fifoOut[31][3];
              muxOutConnector[51] = fifoOut[32][3];
         end
         11: begin
              muxOutConnector[0] = fifoOut[37][15];
              muxOutConnector[1] = fifoOut[38][15];
              muxOutConnector[2] = fifoOut[39][15];
              muxOutConnector[3] = fifoOut[40][15];
              muxOutConnector[4] = fifoOut[41][15];
              muxOutConnector[5] = fifoOut[42][15];
              muxOutConnector[6] = fifoOut[43][15];
              muxOutConnector[7] = fifoOut[44][15];
              muxOutConnector[8] = fifoOut[45][15];
              muxOutConnector[9] = fifoOut[46][15];
              muxOutConnector[10] = fifoOut[47][15];
              muxOutConnector[11] = fifoOut[48][15];
              muxOutConnector[12] = fifoOut[49][15];
              muxOutConnector[13] = fifoOut[50][15];
              muxOutConnector[14] = fifoOut[51][15];
              muxOutConnector[15] = fifoOut[26][14];
              muxOutConnector[16] = fifoOut[27][14];
              muxOutConnector[17] = fifoOut[28][14];
              muxOutConnector[18] = fifoOut[29][14];
              muxOutConnector[19] = fifoOut[30][14];
              muxOutConnector[20] = fifoOut[31][14];
              muxOutConnector[21] = fifoOut[32][14];
              muxOutConnector[22] = fifoOut[33][14];
              muxOutConnector[23] = fifoOut[34][14];
              muxOutConnector[24] = fifoOut[35][14];
              muxOutConnector[25] = fifoOut[36][14];
              muxOutConnector[26] = fifoOut[33][4];
              muxOutConnector[27] = fifoOut[34][4];
              muxOutConnector[28] = fifoOut[35][4];
              muxOutConnector[29] = fifoOut[36][4];
              muxOutConnector[30] = fifoOut[37][4];
              muxOutConnector[31] = fifoOut[38][4];
              muxOutConnector[32] = fifoOut[39][4];
              muxOutConnector[33] = fifoOut[40][4];
              muxOutConnector[34] = fifoOut[41][4];
              muxOutConnector[35] = fifoOut[42][4];
              muxOutConnector[36] = fifoOut[43][4];
              muxOutConnector[37] = fifoOut[44][4];
              muxOutConnector[38] = fifoOut[45][4];
              muxOutConnector[39] = fifoOut[46][4];
              muxOutConnector[40] = fifoOut[47][4];
              muxOutConnector[41] = fifoOut[48][4];
              muxOutConnector[42] = fifoOut[49][4];
              muxOutConnector[43] = fifoOut[50][4];
              muxOutConnector[44] = fifoOut[51][4];
              muxOutConnector[45] = fifoOut[26][3];
              muxOutConnector[46] = fifoOut[27][3];
              muxOutConnector[47] = fifoOut[28][3];
              muxOutConnector[48] = fifoOut[29][3];
              muxOutConnector[49] = fifoOut[30][3];
              muxOutConnector[50] = fifoOut[31][3];
              muxOutConnector[51] = fifoOut[32][3];
         end
         12: begin
              muxOutConnector[0] = fifoOut[37][15];
              muxOutConnector[1] = fifoOut[38][15];
              muxOutConnector[2] = fifoOut[39][15];
              muxOutConnector[3] = fifoOut[40][15];
              muxOutConnector[4] = fifoOut[41][15];
              muxOutConnector[5] = fifoOut[42][15];
              muxOutConnector[6] = fifoOut[43][15];
              muxOutConnector[7] = fifoOut[44][15];
              muxOutConnector[8] = fifoOut[45][15];
              muxOutConnector[9] = fifoOut[46][15];
              muxOutConnector[10] = fifoOut[47][15];
              muxOutConnector[11] = fifoOut[48][15];
              muxOutConnector[12] = fifoOut[49][15];
              muxOutConnector[13] = fifoOut[50][15];
              muxOutConnector[14] = fifoOut[51][15];
              muxOutConnector[15] = fifoOut[26][14];
              muxOutConnector[16] = fifoOut[27][14];
              muxOutConnector[17] = fifoOut[28][14];
              muxOutConnector[18] = fifoOut[29][14];
              muxOutConnector[19] = fifoOut[30][14];
              muxOutConnector[20] = fifoOut[31][14];
              muxOutConnector[21] = fifoOut[32][14];
              muxOutConnector[22] = fifoOut[33][14];
              muxOutConnector[23] = fifoOut[34][14];
              muxOutConnector[24] = fifoOut[35][14];
              muxOutConnector[25] = fifoOut[36][14];
              muxOutConnector[26] = fifoOut[33][4];
              muxOutConnector[27] = fifoOut[34][4];
              muxOutConnector[28] = fifoOut[35][4];
              muxOutConnector[29] = fifoOut[36][4];
              muxOutConnector[30] = fifoOut[37][4];
              muxOutConnector[31] = fifoOut[38][4];
              muxOutConnector[32] = fifoOut[39][4];
              muxOutConnector[33] = fifoOut[40][4];
              muxOutConnector[34] = fifoOut[41][4];
              muxOutConnector[35] = fifoOut[42][4];
              muxOutConnector[36] = fifoOut[43][4];
              muxOutConnector[37] = fifoOut[44][4];
              muxOutConnector[38] = fifoOut[45][4];
              muxOutConnector[39] = fifoOut[46][4];
              muxOutConnector[40] = fifoOut[47][4];
              muxOutConnector[41] = fifoOut[48][4];
              muxOutConnector[42] = fifoOut[49][4];
              muxOutConnector[43] = fifoOut[50][4];
              muxOutConnector[44] = fifoOut[51][4];
              muxOutConnector[45] = fifoOut[26][3];
              muxOutConnector[46] = fifoOut[27][3];
              muxOutConnector[47] = fifoOut[28][3];
              muxOutConnector[48] = fifoOut[29][3];
              muxOutConnector[49] = fifoOut[30][3];
              muxOutConnector[50] = fifoOut[31][3];
              muxOutConnector[51] = fifoOut[32][3];
         end
         13: begin
              muxOutConnector[0] = fifoOut[37][15];
              muxOutConnector[1] = fifoOut[38][15];
              muxOutConnector[2] = fifoOut[39][15];
              muxOutConnector[3] = fifoOut[40][15];
              muxOutConnector[4] = fifoOut[41][15];
              muxOutConnector[5] = fifoOut[42][15];
              muxOutConnector[6] = fifoOut[43][15];
              muxOutConnector[7] = fifoOut[44][15];
              muxOutConnector[8] = fifoOut[45][15];
              muxOutConnector[9] = fifoOut[46][15];
              muxOutConnector[10] = fifoOut[47][15];
              muxOutConnector[11] = fifoOut[48][15];
              muxOutConnector[12] = fifoOut[49][15];
              muxOutConnector[13] = fifoOut[50][15];
              muxOutConnector[14] = fifoOut[51][15];
              muxOutConnector[15] = fifoOut[26][14];
              muxOutConnector[16] = fifoOut[27][14];
              muxOutConnector[17] = fifoOut[28][14];
              muxOutConnector[18] = fifoOut[29][14];
              muxOutConnector[19] = fifoOut[30][14];
              muxOutConnector[20] = fifoOut[31][14];
              muxOutConnector[21] = fifoOut[32][14];
              muxOutConnector[22] = fifoOut[33][14];
              muxOutConnector[23] = fifoOut[34][14];
              muxOutConnector[24] = fifoOut[35][14];
              muxOutConnector[25] = fifoOut[36][14];
              muxOutConnector[26] = fifoOut[33][4];
              muxOutConnector[27] = fifoOut[34][4];
              muxOutConnector[28] = fifoOut[35][4];
              muxOutConnector[29] = fifoOut[36][4];
              muxOutConnector[30] = fifoOut[37][4];
              muxOutConnector[31] = fifoOut[38][4];
              muxOutConnector[32] = fifoOut[39][4];
              muxOutConnector[33] = fifoOut[40][4];
              muxOutConnector[34] = fifoOut[41][4];
              muxOutConnector[35] = fifoOut[42][4];
              muxOutConnector[36] = fifoOut[43][4];
              muxOutConnector[37] = fifoOut[44][4];
              muxOutConnector[38] = fifoOut[45][4];
              muxOutConnector[39] = fifoOut[46][4];
              muxOutConnector[40] = fifoOut[47][4];
              muxOutConnector[41] = fifoOut[48][4];
              muxOutConnector[42] = fifoOut[49][4];
              muxOutConnector[43] = fifoOut[50][4];
              muxOutConnector[44] = fifoOut[51][4];
              muxOutConnector[45] = fifoOut[26][3];
              muxOutConnector[46] = fifoOut[27][3];
              muxOutConnector[47] = fifoOut[28][3];
              muxOutConnector[48] = fifoOut[29][3];
              muxOutConnector[49] = fifoOut[30][3];
              muxOutConnector[50] = fifoOut[31][3];
              muxOutConnector[51] = fifoOut[32][3];
         end
         14: begin
              muxOutConnector[0] = fifoOut[37][15];
              muxOutConnector[1] = fifoOut[38][15];
              muxOutConnector[2] = fifoOut[39][15];
              muxOutConnector[3] = fifoOut[40][15];
              muxOutConnector[4] = fifoOut[41][15];
              muxOutConnector[5] = fifoOut[42][15];
              muxOutConnector[6] = fifoOut[43][15];
              muxOutConnector[7] = fifoOut[44][15];
              muxOutConnector[8] = fifoOut[45][15];
              muxOutConnector[9] = fifoOut[46][15];
              muxOutConnector[10] = fifoOut[47][15];
              muxOutConnector[11] = fifoOut[48][15];
              muxOutConnector[12] = fifoOut[49][15];
              muxOutConnector[13] = fifoOut[50][15];
              muxOutConnector[14] = fifoOut[51][15];
              muxOutConnector[15] = fifoOut[26][14];
              muxOutConnector[16] = fifoOut[27][14];
              muxOutConnector[17] = fifoOut[28][14];
              muxOutConnector[18] = fifoOut[29][14];
              muxOutConnector[19] = fifoOut[30][14];
              muxOutConnector[20] = fifoOut[31][14];
              muxOutConnector[21] = fifoOut[32][14];
              muxOutConnector[22] = fifoOut[33][14];
              muxOutConnector[23] = fifoOut[34][14];
              muxOutConnector[24] = fifoOut[35][14];
              muxOutConnector[25] = fifoOut[36][14];
              muxOutConnector[26] = fifoOut[0][10];
              muxOutConnector[27] = fifoOut[1][10];
              muxOutConnector[28] = fifoOut[2][10];
              muxOutConnector[29] = fifoOut[3][10];
              muxOutConnector[30] = fifoOut[4][10];
              muxOutConnector[31] = fifoOut[5][10];
              muxOutConnector[32] = fifoOut[6][10];
              muxOutConnector[33] = fifoOut[7][10];
              muxOutConnector[34] = fifoOut[8][10];
              muxOutConnector[35] = fifoOut[9][10];
              muxOutConnector[36] = fifoOut[10][10];
              muxOutConnector[37] = fifoOut[11][10];
              muxOutConnector[38] = fifoOut[12][10];
              muxOutConnector[39] = fifoOut[13][10];
              muxOutConnector[40] = fifoOut[14][10];
              muxOutConnector[41] = fifoOut[15][10];
              muxOutConnector[42] = fifoOut[16][10];
              muxOutConnector[43] = fifoOut[17][10];
              muxOutConnector[44] = fifoOut[18][10];
              muxOutConnector[45] = fifoOut[19][10];
              muxOutConnector[46] = fifoOut[20][10];
              muxOutConnector[47] = fifoOut[21][10];
              muxOutConnector[48] = fifoOut[22][10];
              muxOutConnector[49] = fifoOut[23][10];
              muxOutConnector[50] = fifoOut[24][10];
              muxOutConnector[51] = fifoOut[25][10];
         end
         15: begin
              muxOutConnector[0] = fifoOut[37][15];
              muxOutConnector[1] = fifoOut[38][15];
              muxOutConnector[2] = fifoOut[39][15];
              muxOutConnector[3] = fifoOut[40][15];
              muxOutConnector[4] = fifoOut[41][15];
              muxOutConnector[5] = fifoOut[42][15];
              muxOutConnector[6] = fifoOut[10][4];
              muxOutConnector[7] = fifoOut[11][4];
              muxOutConnector[8] = fifoOut[12][4];
              muxOutConnector[9] = fifoOut[13][4];
              muxOutConnector[10] = fifoOut[14][4];
              muxOutConnector[11] = fifoOut[15][4];
              muxOutConnector[12] = fifoOut[16][4];
              muxOutConnector[13] = fifoOut[17][4];
              muxOutConnector[14] = fifoOut[18][4];
              muxOutConnector[15] = fifoOut[19][4];
              muxOutConnector[16] = fifoOut[20][4];
              muxOutConnector[17] = fifoOut[21][4];
              muxOutConnector[18] = fifoOut[22][4];
              muxOutConnector[19] = fifoOut[23][4];
              muxOutConnector[20] = fifoOut[24][4];
              muxOutConnector[21] = fifoOut[25][4];
              muxOutConnector[22] = fifoOut[0][3];
              muxOutConnector[23] = fifoOut[1][3];
              muxOutConnector[24] = fifoOut[2][3];
              muxOutConnector[25] = fifoOut[3][3];
              muxOutConnector[26] = fifoOut[0][10];
              muxOutConnector[27] = fifoOut[1][10];
              muxOutConnector[28] = fifoOut[2][10];
              muxOutConnector[29] = fifoOut[3][10];
              muxOutConnector[30] = fifoOut[4][10];
              muxOutConnector[31] = fifoOut[5][10];
              muxOutConnector[32] = fifoOut[6][10];
              muxOutConnector[33] = fifoOut[7][10];
              muxOutConnector[34] = fifoOut[8][10];
              muxOutConnector[35] = fifoOut[9][10];
              muxOutConnector[36] = fifoOut[10][10];
              muxOutConnector[37] = fifoOut[11][10];
              muxOutConnector[38] = fifoOut[12][10];
              muxOutConnector[39] = fifoOut[13][10];
              muxOutConnector[40] = fifoOut[14][10];
              muxOutConnector[41] = fifoOut[15][10];
              muxOutConnector[42] = fifoOut[16][10];
              muxOutConnector[43] = fifoOut[17][10];
              muxOutConnector[44] = fifoOut[18][10];
              muxOutConnector[45] = fifoOut[19][10];
              muxOutConnector[46] = fifoOut[20][10];
              muxOutConnector[47] = fifoOut[21][10];
              muxOutConnector[48] = fifoOut[22][10];
              muxOutConnector[49] = fifoOut[23][10];
              muxOutConnector[50] = fifoOut[24][10];
              muxOutConnector[51] = fifoOut[25][10];
         end
         16: begin
              muxOutConnector[0] = fifoOut[4][4];
              muxOutConnector[1] = fifoOut[5][4];
              muxOutConnector[2] = fifoOut[6][4];
              muxOutConnector[3] = fifoOut[7][4];
              muxOutConnector[4] = fifoOut[8][4];
              muxOutConnector[5] = fifoOut[9][4];
              muxOutConnector[6] = fifoOut[10][4];
              muxOutConnector[7] = fifoOut[11][4];
              muxOutConnector[8] = fifoOut[12][4];
              muxOutConnector[9] = fifoOut[13][4];
              muxOutConnector[10] = fifoOut[14][4];
              muxOutConnector[11] = fifoOut[15][4];
              muxOutConnector[12] = fifoOut[16][4];
              muxOutConnector[13] = fifoOut[17][4];
              muxOutConnector[14] = fifoOut[18][4];
              muxOutConnector[15] = fifoOut[19][4];
              muxOutConnector[16] = fifoOut[20][4];
              muxOutConnector[17] = fifoOut[21][4];
              muxOutConnector[18] = fifoOut[22][4];
              muxOutConnector[19] = fifoOut[23][4];
              muxOutConnector[20] = fifoOut[24][4];
              muxOutConnector[21] = fifoOut[25][4];
              muxOutConnector[22] = fifoOut[0][3];
              muxOutConnector[23] = fifoOut[1][3];
              muxOutConnector[24] = fifoOut[2][3];
              muxOutConnector[25] = fifoOut[3][3];
              muxOutConnector[26] = fifoOut[0][10];
              muxOutConnector[27] = fifoOut[1][10];
              muxOutConnector[28] = fifoOut[2][10];
              muxOutConnector[29] = fifoOut[3][10];
              muxOutConnector[30] = fifoOut[4][10];
              muxOutConnector[31] = fifoOut[5][10];
              muxOutConnector[32] = fifoOut[6][10];
              muxOutConnector[33] = fifoOut[7][10];
              muxOutConnector[34] = fifoOut[8][10];
              muxOutConnector[35] = fifoOut[9][10];
              muxOutConnector[36] = fifoOut[10][10];
              muxOutConnector[37] = fifoOut[11][10];
              muxOutConnector[38] = fifoOut[12][10];
              muxOutConnector[39] = fifoOut[13][10];
              muxOutConnector[40] = fifoOut[14][10];
              muxOutConnector[41] = fifoOut[15][10];
              muxOutConnector[42] = fifoOut[16][10];
              muxOutConnector[43] = fifoOut[17][10];
              muxOutConnector[44] = fifoOut[18][10];
              muxOutConnector[45] = fifoOut[19][10];
              muxOutConnector[46] = fifoOut[20][10];
              muxOutConnector[47] = fifoOut[21][10];
              muxOutConnector[48] = fifoOut[22][10];
              muxOutConnector[49] = fifoOut[23][10];
              muxOutConnector[50] = fifoOut[24][10];
              muxOutConnector[51] = fifoOut[25][10];
         end
         17: begin
              muxOutConnector[0] = fifoOut[4][4];
              muxOutConnector[1] = fifoOut[5][4];
              muxOutConnector[2] = fifoOut[6][4];
              muxOutConnector[3] = fifoOut[7][4];
              muxOutConnector[4] = fifoOut[8][4];
              muxOutConnector[5] = fifoOut[9][4];
              muxOutConnector[6] = fifoOut[10][4];
              muxOutConnector[7] = fifoOut[11][4];
              muxOutConnector[8] = fifoOut[12][4];
              muxOutConnector[9] = fifoOut[13][4];
              muxOutConnector[10] = fifoOut[14][4];
              muxOutConnector[11] = fifoOut[15][4];
              muxOutConnector[12] = fifoOut[16][4];
              muxOutConnector[13] = fifoOut[17][4];
              muxOutConnector[14] = fifoOut[18][4];
              muxOutConnector[15] = fifoOut[19][4];
              muxOutConnector[16] = fifoOut[20][4];
              muxOutConnector[17] = fifoOut[21][4];
              muxOutConnector[18] = fifoOut[22][4];
              muxOutConnector[19] = fifoOut[23][4];
              muxOutConnector[20] = fifoOut[24][4];
              muxOutConnector[21] = fifoOut[25][4];
              muxOutConnector[22] = fifoOut[0][3];
              muxOutConnector[23] = fifoOut[1][3];
              muxOutConnector[24] = fifoOut[2][3];
              muxOutConnector[25] = fifoOut[3][3];
              muxOutConnector[26] = fifoOut[0][10];
              muxOutConnector[27] = fifoOut[1][10];
              muxOutConnector[28] = fifoOut[2][10];
              muxOutConnector[29] = fifoOut[3][10];
              muxOutConnector[30] = fifoOut[4][10];
              muxOutConnector[31] = fifoOut[5][10];
              muxOutConnector[32] = fifoOut[6][10];
              muxOutConnector[33] = fifoOut[7][10];
              muxOutConnector[34] = fifoOut[8][10];
              muxOutConnector[35] = fifoOut[9][10];
              muxOutConnector[36] = fifoOut[10][10];
              muxOutConnector[37] = fifoOut[11][10];
              muxOutConnector[38] = fifoOut[12][10];
              muxOutConnector[39] = fifoOut[13][10];
              muxOutConnector[40] = fifoOut[14][10];
              muxOutConnector[41] = fifoOut[15][10];
              muxOutConnector[42] = fifoOut[16][10];
              muxOutConnector[43] = fifoOut[17][10];
              muxOutConnector[44] = fifoOut[18][10];
              muxOutConnector[45] = fifoOut[19][10];
              muxOutConnector[46] = fifoOut[20][10];
              muxOutConnector[47] = fifoOut[21][10];
              muxOutConnector[48] = fifoOut[22][10];
              muxOutConnector[49] = fifoOut[23][10];
              muxOutConnector[50] = fifoOut[24][10];
              muxOutConnector[51] = fifoOut[25][10];
         end
         18: begin
              muxOutConnector[0] = fifoOut[4][4];
              muxOutConnector[1] = fifoOut[5][4];
              muxOutConnector[2] = fifoOut[6][4];
              muxOutConnector[3] = fifoOut[7][4];
              muxOutConnector[4] = fifoOut[8][4];
              muxOutConnector[5] = fifoOut[9][4];
              muxOutConnector[6] = fifoOut[10][4];
              muxOutConnector[7] = fifoOut[11][4];
              muxOutConnector[8] = fifoOut[12][4];
              muxOutConnector[9] = fifoOut[13][4];
              muxOutConnector[10] = fifoOut[14][4];
              muxOutConnector[11] = fifoOut[15][4];
              muxOutConnector[12] = fifoOut[16][4];
              muxOutConnector[13] = fifoOut[17][4];
              muxOutConnector[14] = fifoOut[18][4];
              muxOutConnector[15] = fifoOut[19][4];
              muxOutConnector[16] = fifoOut[20][4];
              muxOutConnector[17] = fifoOut[21][4];
              muxOutConnector[18] = fifoOut[22][4];
              muxOutConnector[19] = fifoOut[23][4];
              muxOutConnector[20] = fifoOut[24][4];
              muxOutConnector[21] = fifoOut[25][4];
              muxOutConnector[22] = fifoOut[0][3];
              muxOutConnector[23] = fifoOut[1][3];
              muxOutConnector[24] = fifoOut[2][3];
              muxOutConnector[25] = fifoOut[3][3];
              muxOutConnector[26] = fifoOut[0][10];
              muxOutConnector[27] = fifoOut[1][10];
              muxOutConnector[28] = fifoOut[2][10];
              muxOutConnector[29] = fifoOut[3][10];
              muxOutConnector[30] = fifoOut[4][10];
              muxOutConnector[31] = fifoOut[5][10];
              muxOutConnector[32] = fifoOut[6][10];
              muxOutConnector[33] = fifoOut[7][10];
              muxOutConnector[34] = fifoOut[8][10];
              muxOutConnector[35] = fifoOut[9][10];
              muxOutConnector[36] = fifoOut[10][10];
              muxOutConnector[37] = fifoOut[11][10];
              muxOutConnector[38] = fifoOut[12][10];
              muxOutConnector[39] = fifoOut[13][10];
              muxOutConnector[40] = fifoOut[14][10];
              muxOutConnector[41] = fifoOut[15][10];
              muxOutConnector[42] = fifoOut[16][10];
              muxOutConnector[43] = fifoOut[17][10];
              muxOutConnector[44] = fifoOut[18][10];
              muxOutConnector[45] = fifoOut[19][10];
              muxOutConnector[46] = fifoOut[20][10];
              muxOutConnector[47] = fifoOut[21][10];
              muxOutConnector[48] = fifoOut[22][10];
              muxOutConnector[49] = fifoOut[23][10];
              muxOutConnector[50] = fifoOut[24][10];
              muxOutConnector[51] = fifoOut[25][10];
         end
         19: begin
              muxOutConnector[0] = fifoOut[4][4];
              muxOutConnector[1] = fifoOut[5][4];
              muxOutConnector[2] = fifoOut[6][4];
              muxOutConnector[3] = fifoOut[7][4];
              muxOutConnector[4] = fifoOut[8][4];
              muxOutConnector[5] = fifoOut[9][4];
              muxOutConnector[6] = fifoOut[10][4];
              muxOutConnector[7] = fifoOut[11][4];
              muxOutConnector[8] = fifoOut[12][4];
              muxOutConnector[9] = fifoOut[13][4];
              muxOutConnector[10] = fifoOut[14][4];
              muxOutConnector[11] = fifoOut[15][4];
              muxOutConnector[12] = fifoOut[16][4];
              muxOutConnector[13] = fifoOut[17][4];
              muxOutConnector[14] = fifoOut[18][4];
              muxOutConnector[15] = fifoOut[19][4];
              muxOutConnector[16] = fifoOut[20][4];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[0][10];
              muxOutConnector[27] = fifoOut[1][10];
              muxOutConnector[28] = fifoOut[2][10];
              muxOutConnector[29] = fifoOut[3][10];
              muxOutConnector[30] = fifoOut[4][10];
              muxOutConnector[31] = fifoOut[5][10];
              muxOutConnector[32] = fifoOut[6][10];
              muxOutConnector[33] = fifoOut[7][10];
              muxOutConnector[34] = fifoOut[8][10];
              muxOutConnector[35] = fifoOut[9][10];
              muxOutConnector[36] = fifoOut[10][10];
              muxOutConnector[37] = fifoOut[11][10];
              muxOutConnector[38] = fifoOut[12][10];
              muxOutConnector[39] = fifoOut[13][10];
              muxOutConnector[40] = fifoOut[14][10];
              muxOutConnector[41] = fifoOut[15][10];
              muxOutConnector[42] = fifoOut[16][10];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
         end
         default: begin
               for(i=0;i<muxOutSymbols;i=i+1)begin
                muxOutConnector[i] = 0;
              end
         end
//hgjhgbuiguigbigbgbgbui
         endcase
    end
endcase
             end
        endmodule