`timescale 1ns / 1ps
/////////////////////////////////////////////////
//script: circulant_shiftregAlign.m
/////////////////////////////////////////////////
module writeselector_inputintf(wr_en_vec,wr_address_vec,cyclecount,wr_en);
parameter ADDRESSWIDTH = 5;
//Non-configurable
parameter Nb = 16;//16*511=8176 codeword

parameter CYCLECOUNTWIDTH = 8;//maxcycles=(8160+32)/32)=256, width=ceil(log2(256))=8

output reg[Nb-1:0] wr_en_vec;
output [(Nb*ADDRESSWIDTH)-1:0] wr_address_vec;
input[(CYCLECOUNTWIDTH)-1:0] cyclecount;
input wr_en;

reg[(ADDRESSWIDTH)-1:0] wr_address[Nb-1:0];
genvar i;
generate
    for (i=0;i<Nb;i=i+1)begin:nb_loop
        assign wr_address_vec[ ((i+1)*ADDRESSWIDTH)-1:i*ADDRESSWIDTH]=wr_address[i];
    end
endgenerate

always@(*) begin
  case(cyclecount)
   1: begin
         wr_en_vec[0]=1;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   2: begin
         wr_en_vec[0]=1;
         wr_address[0]=1;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   3: begin
         wr_en_vec[0]=1;
         wr_address[0]=2;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   4: begin
         wr_en_vec[0]=1;
         wr_address[0]=3;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   5: begin
         wr_en_vec[0]=1;
         wr_address[0]=4;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   6: begin
         wr_en_vec[0]=1;
         wr_address[0]=5;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   7: begin
         wr_en_vec[0]=1;
         wr_address[0]=6;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   8: begin
         wr_en_vec[0]=1;
         wr_address[0]=7;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   9: begin
         wr_en_vec[0]=1;
         wr_address[0]=8;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   10: begin
         wr_en_vec[0]=1;
         wr_address[0]=9;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   11: begin
         wr_en_vec[0]=1;
         wr_address[0]=10;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   12: begin
         wr_en_vec[0]=1;
         wr_address[0]=11;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   13: begin
         wr_en_vec[0]=1;
         wr_address[0]=12;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   14: begin
         wr_en_vec[0]=1;
         wr_address[0]=13;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   15: begin
         wr_en_vec[0]=1;
         wr_address[0]=14;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   16: begin
         wr_en_vec[0]=1;
         wr_address[0]=15;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   17: begin
         wr_en_vec[1]=1;
         wr_address[1]=0;
         wr_en_vec[0]=1;
         wr_address[0]=16;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   18: begin
         wr_en_vec[1]=1;
         wr_address[1]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   19: begin
         wr_en_vec[1]=1;
         wr_address[1]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   20: begin
         wr_en_vec[1]=1;
         wr_address[1]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   21: begin
         wr_en_vec[1]=1;
         wr_address[1]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   22: begin
         wr_en_vec[1]=1;
         wr_address[1]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   23: begin
         wr_en_vec[1]=1;
         wr_address[1]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   24: begin
         wr_en_vec[1]=1;
         wr_address[1]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   25: begin
         wr_en_vec[1]=1;
         wr_address[1]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   26: begin
         wr_en_vec[1]=1;
         wr_address[1]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   27: begin
         wr_en_vec[1]=1;
         wr_address[1]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   28: begin
         wr_en_vec[1]=1;
         wr_address[1]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   29: begin
         wr_en_vec[1]=1;
         wr_address[1]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   30: begin
         wr_en_vec[1]=1;
         wr_address[1]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   31: begin
         wr_en_vec[1]=1;
         wr_address[1]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   32: begin
         wr_en_vec[1]=1;
         wr_address[1]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   33: begin
         wr_en_vec[2]=1;
         wr_address[2]=0;
         wr_en_vec[1]=1;
         wr_address[1]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   34: begin
         wr_en_vec[2]=1;
         wr_address[2]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   35: begin
         wr_en_vec[2]=1;
         wr_address[2]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   36: begin
         wr_en_vec[2]=1;
         wr_address[2]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   37: begin
         wr_en_vec[2]=1;
         wr_address[2]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   38: begin
         wr_en_vec[2]=1;
         wr_address[2]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   39: begin
         wr_en_vec[2]=1;
         wr_address[2]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   40: begin
         wr_en_vec[2]=1;
         wr_address[2]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   41: begin
         wr_en_vec[2]=1;
         wr_address[2]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   42: begin
         wr_en_vec[2]=1;
         wr_address[2]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   43: begin
         wr_en_vec[2]=1;
         wr_address[2]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   44: begin
         wr_en_vec[2]=1;
         wr_address[2]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   45: begin
         wr_en_vec[2]=1;
         wr_address[2]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   46: begin
         wr_en_vec[2]=1;
         wr_address[2]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   47: begin
         wr_en_vec[2]=1;
         wr_address[2]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   48: begin
         wr_en_vec[2]=1;
         wr_address[2]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   49: begin
         wr_en_vec[3]=1;
         wr_address[3]=0;
         wr_en_vec[2]=1;
         wr_address[2]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   50: begin
         wr_en_vec[3]=1;
         wr_address[3]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   51: begin
         wr_en_vec[3]=1;
         wr_address[3]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   52: begin
         wr_en_vec[3]=1;
         wr_address[3]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   53: begin
         wr_en_vec[3]=1;
         wr_address[3]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   54: begin
         wr_en_vec[3]=1;
         wr_address[3]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   55: begin
         wr_en_vec[3]=1;
         wr_address[3]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   56: begin
         wr_en_vec[3]=1;
         wr_address[3]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   57: begin
         wr_en_vec[3]=1;
         wr_address[3]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   58: begin
         wr_en_vec[3]=1;
         wr_address[3]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   59: begin
         wr_en_vec[3]=1;
         wr_address[3]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   60: begin
         wr_en_vec[3]=1;
         wr_address[3]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   61: begin
         wr_en_vec[3]=1;
         wr_address[3]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   62: begin
         wr_en_vec[3]=1;
         wr_address[3]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   63: begin
         wr_en_vec[3]=1;
         wr_address[3]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   64: begin
         wr_en_vec[3]=1;
         wr_address[3]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   65: begin
         wr_en_vec[4]=1;
         wr_address[4]=0;
         wr_en_vec[3]=1;
         wr_address[3]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   66: begin
         wr_en_vec[4]=1;
         wr_address[4]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   67: begin
         wr_en_vec[4]=1;
         wr_address[4]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   68: begin
         wr_en_vec[4]=1;
         wr_address[4]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   69: begin
         wr_en_vec[4]=1;
         wr_address[4]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   70: begin
         wr_en_vec[4]=1;
         wr_address[4]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   71: begin
         wr_en_vec[4]=1;
         wr_address[4]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   72: begin
         wr_en_vec[4]=1;
         wr_address[4]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   73: begin
         wr_en_vec[4]=1;
         wr_address[4]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   74: begin
         wr_en_vec[4]=1;
         wr_address[4]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   75: begin
         wr_en_vec[4]=1;
         wr_address[4]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   76: begin
         wr_en_vec[4]=1;
         wr_address[4]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   77: begin
         wr_en_vec[4]=1;
         wr_address[4]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   78: begin
         wr_en_vec[4]=1;
         wr_address[4]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   79: begin
         wr_en_vec[4]=1;
         wr_address[4]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   80: begin
         wr_en_vec[4]=1;
         wr_address[4]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   81: begin
         wr_en_vec[5]=1;
         wr_address[5]=0;
         wr_en_vec[4]=1;
         wr_address[4]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   82: begin
         wr_en_vec[5]=1;
         wr_address[5]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   83: begin
         wr_en_vec[5]=1;
         wr_address[5]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   84: begin
         wr_en_vec[5]=1;
         wr_address[5]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   85: begin
         wr_en_vec[5]=1;
         wr_address[5]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   86: begin
         wr_en_vec[5]=1;
         wr_address[5]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   87: begin
         wr_en_vec[5]=1;
         wr_address[5]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   88: begin
         wr_en_vec[5]=1;
         wr_address[5]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   89: begin
         wr_en_vec[5]=1;
         wr_address[5]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   90: begin
         wr_en_vec[5]=1;
         wr_address[5]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   91: begin
         wr_en_vec[5]=1;
         wr_address[5]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   92: begin
         wr_en_vec[5]=1;
         wr_address[5]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   93: begin
         wr_en_vec[5]=1;
         wr_address[5]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   94: begin
         wr_en_vec[5]=1;
         wr_address[5]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   95: begin
         wr_en_vec[5]=1;
         wr_address[5]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   96: begin
         wr_en_vec[5]=1;
         wr_address[5]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   97: begin
         wr_en_vec[6]=1;
         wr_address[6]=0;
         wr_en_vec[5]=1;
         wr_address[5]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   98: begin
         wr_en_vec[6]=1;
         wr_address[6]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   99: begin
         wr_en_vec[6]=1;
         wr_address[6]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   100: begin
         wr_en_vec[6]=1;
         wr_address[6]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   101: begin
         wr_en_vec[6]=1;
         wr_address[6]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   102: begin
         wr_en_vec[6]=1;
         wr_address[6]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   103: begin
         wr_en_vec[6]=1;
         wr_address[6]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   104: begin
         wr_en_vec[6]=1;
         wr_address[6]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   105: begin
         wr_en_vec[6]=1;
         wr_address[6]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   106: begin
         wr_en_vec[6]=1;
         wr_address[6]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   107: begin
         wr_en_vec[6]=1;
         wr_address[6]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   108: begin
         wr_en_vec[6]=1;
         wr_address[6]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   109: begin
         wr_en_vec[6]=1;
         wr_address[6]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   110: begin
         wr_en_vec[6]=1;
         wr_address[6]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   111: begin
         wr_en_vec[6]=1;
         wr_address[6]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   112: begin
         wr_en_vec[6]=1;
         wr_address[6]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   113: begin
         wr_en_vec[7]=1;
         wr_address[7]=0;
         wr_en_vec[6]=1;
         wr_address[6]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   114: begin
         wr_en_vec[7]=1;
         wr_address[7]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   115: begin
         wr_en_vec[7]=1;
         wr_address[7]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   116: begin
         wr_en_vec[7]=1;
         wr_address[7]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   117: begin
         wr_en_vec[7]=1;
         wr_address[7]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   118: begin
         wr_en_vec[7]=1;
         wr_address[7]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   119: begin
         wr_en_vec[7]=1;
         wr_address[7]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   120: begin
         wr_en_vec[7]=1;
         wr_address[7]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   121: begin
         wr_en_vec[7]=1;
         wr_address[7]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   122: begin
         wr_en_vec[7]=1;
         wr_address[7]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   123: begin
         wr_en_vec[7]=1;
         wr_address[7]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   124: begin
         wr_en_vec[7]=1;
         wr_address[7]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   125: begin
         wr_en_vec[7]=1;
         wr_address[7]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   126: begin
         wr_en_vec[7]=1;
         wr_address[7]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   127: begin
         wr_en_vec[7]=1;
         wr_address[7]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   128: begin
         wr_en_vec[7]=1;
         wr_address[7]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   129: begin
         wr_en_vec[8]=1;
         wr_address[8]=0;
         wr_en_vec[7]=1;
         wr_address[7]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   130: begin
         wr_en_vec[8]=1;
         wr_address[8]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   131: begin
         wr_en_vec[8]=1;
         wr_address[8]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   132: begin
         wr_en_vec[8]=1;
         wr_address[8]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   133: begin
         wr_en_vec[8]=1;
         wr_address[8]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   134: begin
         wr_en_vec[8]=1;
         wr_address[8]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   135: begin
         wr_en_vec[8]=1;
         wr_address[8]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   136: begin
         wr_en_vec[8]=1;
         wr_address[8]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   137: begin
         wr_en_vec[8]=1;
         wr_address[8]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   138: begin
         wr_en_vec[8]=1;
         wr_address[8]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   139: begin
         wr_en_vec[8]=1;
         wr_address[8]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   140: begin
         wr_en_vec[8]=1;
         wr_address[8]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   141: begin
         wr_en_vec[8]=1;
         wr_address[8]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   142: begin
         wr_en_vec[8]=1;
         wr_address[8]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   143: begin
         wr_en_vec[8]=1;
         wr_address[8]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   144: begin
         wr_en_vec[8]=1;
         wr_address[8]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   145: begin
         wr_en_vec[9]=1;
         wr_address[9]=0;
         wr_en_vec[8]=1;
         wr_address[8]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   146: begin
         wr_en_vec[9]=1;
         wr_address[9]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   147: begin
         wr_en_vec[9]=1;
         wr_address[9]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   148: begin
         wr_en_vec[9]=1;
         wr_address[9]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   149: begin
         wr_en_vec[9]=1;
         wr_address[9]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   150: begin
         wr_en_vec[9]=1;
         wr_address[9]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   151: begin
         wr_en_vec[9]=1;
         wr_address[9]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   152: begin
         wr_en_vec[9]=1;
         wr_address[9]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   153: begin
         wr_en_vec[9]=1;
         wr_address[9]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   154: begin
         wr_en_vec[9]=1;
         wr_address[9]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   155: begin
         wr_en_vec[9]=1;
         wr_address[9]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   156: begin
         wr_en_vec[9]=1;
         wr_address[9]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   157: begin
         wr_en_vec[9]=1;
         wr_address[9]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   158: begin
         wr_en_vec[9]=1;
         wr_address[9]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   159: begin
         wr_en_vec[9]=1;
         wr_address[9]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   160: begin
         wr_en_vec[9]=1;
         wr_address[9]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   161: begin
         wr_en_vec[10]=1;
         wr_address[10]=0;
         wr_en_vec[9]=1;
         wr_address[9]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   162: begin
         wr_en_vec[10]=1;
         wr_address[10]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   163: begin
         wr_en_vec[10]=1;
         wr_address[10]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   164: begin
         wr_en_vec[10]=1;
         wr_address[10]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   165: begin
         wr_en_vec[10]=1;
         wr_address[10]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   166: begin
         wr_en_vec[10]=1;
         wr_address[10]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   167: begin
         wr_en_vec[10]=1;
         wr_address[10]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   168: begin
         wr_en_vec[10]=1;
         wr_address[10]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   169: begin
         wr_en_vec[10]=1;
         wr_address[10]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   170: begin
         wr_en_vec[10]=1;
         wr_address[10]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   171: begin
         wr_en_vec[10]=1;
         wr_address[10]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   172: begin
         wr_en_vec[10]=1;
         wr_address[10]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   173: begin
         wr_en_vec[10]=1;
         wr_address[10]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   174: begin
         wr_en_vec[10]=1;
         wr_address[10]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   175: begin
         wr_en_vec[10]=1;
         wr_address[10]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   176: begin
         wr_en_vec[10]=1;
         wr_address[10]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   177: begin
         wr_en_vec[11]=1;
         wr_address[11]=0;
         wr_en_vec[10]=1;
         wr_address[10]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   178: begin
         wr_en_vec[11]=1;
         wr_address[11]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   179: begin
         wr_en_vec[11]=1;
         wr_address[11]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   180: begin
         wr_en_vec[11]=1;
         wr_address[11]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   181: begin
         wr_en_vec[11]=1;
         wr_address[11]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   182: begin
         wr_en_vec[11]=1;
         wr_address[11]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   183: begin
         wr_en_vec[11]=1;
         wr_address[11]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   184: begin
         wr_en_vec[11]=1;
         wr_address[11]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   185: begin
         wr_en_vec[11]=1;
         wr_address[11]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   186: begin
         wr_en_vec[11]=1;
         wr_address[11]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   187: begin
         wr_en_vec[11]=1;
         wr_address[11]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   188: begin
         wr_en_vec[11]=1;
         wr_address[11]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   189: begin
         wr_en_vec[11]=1;
         wr_address[11]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   190: begin
         wr_en_vec[11]=1;
         wr_address[11]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   191: begin
         wr_en_vec[11]=1;
         wr_address[11]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   192: begin
         wr_en_vec[11]=1;
         wr_address[11]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   193: begin
         wr_en_vec[12]=1;
         wr_address[12]=0;
         wr_en_vec[11]=1;
         wr_address[11]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   194: begin
         wr_en_vec[12]=1;
         wr_address[12]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   195: begin
         wr_en_vec[12]=1;
         wr_address[12]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   196: begin
         wr_en_vec[12]=1;
         wr_address[12]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   197: begin
         wr_en_vec[12]=1;
         wr_address[12]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   198: begin
         wr_en_vec[12]=1;
         wr_address[12]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   199: begin
         wr_en_vec[12]=1;
         wr_address[12]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   200: begin
         wr_en_vec[12]=1;
         wr_address[12]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   201: begin
         wr_en_vec[12]=1;
         wr_address[12]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   202: begin
         wr_en_vec[12]=1;
         wr_address[12]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   203: begin
         wr_en_vec[12]=1;
         wr_address[12]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   204: begin
         wr_en_vec[12]=1;
         wr_address[12]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   205: begin
         wr_en_vec[12]=1;
         wr_address[12]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   206: begin
         wr_en_vec[12]=1;
         wr_address[12]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   207: begin
         wr_en_vec[12]=1;
         wr_address[12]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   208: begin
         wr_en_vec[12]=1;
         wr_address[12]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   209: begin
         wr_en_vec[13]=1;
         wr_address[13]=0;
         wr_en_vec[12]=1;
         wr_address[12]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   210: begin
         wr_en_vec[13]=1;
         wr_address[13]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   211: begin
         wr_en_vec[13]=1;
         wr_address[13]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   212: begin
         wr_en_vec[13]=1;
         wr_address[13]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   213: begin
         wr_en_vec[13]=1;
         wr_address[13]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   214: begin
         wr_en_vec[13]=1;
         wr_address[13]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   215: begin
         wr_en_vec[13]=1;
         wr_address[13]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   216: begin
         wr_en_vec[13]=1;
         wr_address[13]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   217: begin
         wr_en_vec[13]=1;
         wr_address[13]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   218: begin
         wr_en_vec[13]=1;
         wr_address[13]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   219: begin
         wr_en_vec[13]=1;
         wr_address[13]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   220: begin
         wr_en_vec[13]=1;
         wr_address[13]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   221: begin
         wr_en_vec[13]=1;
         wr_address[13]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   222: begin
         wr_en_vec[13]=1;
         wr_address[13]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   223: begin
         wr_en_vec[13]=1;
         wr_address[13]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   224: begin
         wr_en_vec[13]=1;
         wr_address[13]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   225: begin
         wr_en_vec[14]=1;
         wr_address[14]=0;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   226: begin
         wr_en_vec[14]=1;
         wr_address[14]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   227: begin
         wr_en_vec[14]=1;
         wr_address[14]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   228: begin
         wr_en_vec[14]=1;
         wr_address[14]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   229: begin
         wr_en_vec[14]=1;
         wr_address[14]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   230: begin
         wr_en_vec[14]=1;
         wr_address[14]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   231: begin
         wr_en_vec[14]=1;
         wr_address[14]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   232: begin
         wr_en_vec[14]=1;
         wr_address[14]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   233: begin
         wr_en_vec[14]=1;
         wr_address[14]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   234: begin
         wr_en_vec[14]=1;
         wr_address[14]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   235: begin
         wr_en_vec[14]=1;
         wr_address[14]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   236: begin
         wr_en_vec[14]=1;
         wr_address[14]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   237: begin
         wr_en_vec[14]=1;
         wr_address[14]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   238: begin
         wr_en_vec[14]=1;
         wr_address[14]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   239: begin
         wr_en_vec[14]=1;
         wr_address[14]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   240: begin
         wr_en_vec[15]=1;
         wr_address[15]=0;
         wr_en_vec[14]=1;
         wr_address[14]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
       end
   241: begin
         wr_en_vec[15]=1;
         wr_address[15]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   242: begin
         wr_en_vec[15]=1;
         wr_address[15]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   243: begin
         wr_en_vec[15]=1;
         wr_address[15]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   244: begin
         wr_en_vec[15]=1;
         wr_address[15]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   245: begin
         wr_en_vec[15]=1;
         wr_address[15]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   246: begin
         wr_en_vec[15]=1;
         wr_address[15]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   247: begin
         wr_en_vec[15]=1;
         wr_address[15]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   248: begin
         wr_en_vec[15]=1;
         wr_address[15]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   249: begin
         wr_en_vec[15]=1;
         wr_address[15]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   250: begin
         wr_en_vec[15]=1;
         wr_address[15]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   251: begin
         wr_en_vec[15]=1;
         wr_address[15]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   252: begin
         wr_en_vec[15]=1;
         wr_address[15]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   253: begin
         wr_en_vec[15]=1;
         wr_address[15]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   254: begin
         wr_en_vec[15]=1;
         wr_address[15]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   255: begin
         wr_en_vec[15]=1;
         wr_address[15]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   256: begin
         wr_en_vec[15]=1;
         wr_address[15]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   default: begin
              wr_en_vec[0]=0;
              wr_address[0]=0;
              wr_en_vec[1]=0;
              wr_address[1]=0;
              wr_en_vec[2]=0;
              wr_address[2]=0;
              wr_en_vec[3]=0;
              wr_address[3]=0;
              wr_en_vec[4]=0;
              wr_address[4]=0;
              wr_en_vec[5]=0;
              wr_address[5]=0;
              wr_en_vec[6]=0;
              wr_address[6]=0;
              wr_en_vec[7]=0;
              wr_address[7]=0;
              wr_en_vec[8]=0;
              wr_address[8]=0;
              wr_en_vec[9]=0;
              wr_address[9]=0;
              wr_en_vec[10]=0;
              wr_address[10]=0;
              wr_en_vec[11]=0;
              wr_address[11]=0;
              wr_en_vec[12]=0;
              wr_address[12]=0;
              wr_en_vec[13]=0;
              wr_address[13]=0;
              wr_en_vec[14]=0;
              wr_address[14]=0;
              wr_en_vec[15]=0;
              wr_address[15]=0;
            //first 64 ASM symbols of 0th cycle is skipped using this default case.
            end
  endcase
end

endmodule
