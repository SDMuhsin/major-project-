`timescale 1ns / 1ps
module LMem1To0_511_circ0_ys_yu_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        wr_en,
        feedback_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 15;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input [ADDRESSWIDTH-1:0]unloadAddress;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

input feedback_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        if(feedback_en) begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= fifoOut[i][c-1];
         end
        end
        else begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= ly0InConnector[i];
         end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
       0: begin
              unloadMuxOut[0] = fifoOut[22][4][w-1];
              unloadMuxOut[1] = fifoOut[23][4][w-1];
              unloadMuxOut[2] = fifoOut[24][4][w-1];
              unloadMuxOut[3] = fifoOut[25][4][w-1];
              unloadMuxOut[4] = fifoOut[0][3][w-1];
              unloadMuxOut[5] = fifoOut[1][3][w-1];
              unloadMuxOut[6] = fifoOut[2][3][w-1];
              unloadMuxOut[7] = fifoOut[3][3][w-1];
              unloadMuxOut[8] = fifoOut[4][3][w-1];
              unloadMuxOut[9] = fifoOut[5][3][w-1];
              unloadMuxOut[10] = fifoOut[6][3][w-1];
              unloadMuxOut[11] = fifoOut[7][3][w-1];
              unloadMuxOut[12] = fifoOut[8][3][w-1];
              unloadMuxOut[13] = fifoOut[9][3][w-1];
              unloadMuxOut[14] = fifoOut[10][3][w-1];
              unloadMuxOut[15] = fifoOut[11][3][w-1];
              unloadMuxOut[16] = fifoOut[12][3][w-1];
              unloadMuxOut[17] = fifoOut[13][3][w-1];
              unloadMuxOut[18] = fifoOut[14][3][w-1];
              unloadMuxOut[19] = fifoOut[15][3][w-1];
              unloadMuxOut[20] = fifoOut[16][3][w-1];
              unloadMuxOut[21] = fifoOut[17][3][w-1];
              unloadMuxOut[22] = fifoOut[18][3][w-1];
              unloadMuxOut[23] = fifoOut[19][3][w-1];
              unloadMuxOut[24] = fifoOut[20][3][w-1];
              unloadMuxOut[25] = fifoOut[21][3][w-1];
              unloadMuxOut[26] = fifoOut[22][3][w-1];
              unloadMuxOut[27] = fifoOut[23][3][w-1];
              unloadMuxOut[28] = fifoOut[24][3][w-1];
              unloadMuxOut[29] = fifoOut[25][3][w-1];
              unloadMuxOut[30] = fifoOut[0][2][w-1];
              unloadMuxOut[31] = fifoOut[1][2][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[2][2][w-1];
              unloadMuxOut[1] = fifoOut[3][2][w-1];
              unloadMuxOut[2] = fifoOut[4][2][w-1];
              unloadMuxOut[3] = fifoOut[5][2][w-1];
              unloadMuxOut[4] = fifoOut[6][2][w-1];
              unloadMuxOut[5] = fifoOut[7][2][w-1];
              unloadMuxOut[6] = fifoOut[8][2][w-1];
              unloadMuxOut[7] = fifoOut[9][2][w-1];
              unloadMuxOut[8] = fifoOut[10][2][w-1];
              unloadMuxOut[9] = fifoOut[11][2][w-1];
              unloadMuxOut[10] = fifoOut[12][2][w-1];
              unloadMuxOut[11] = fifoOut[13][2][w-1];
              unloadMuxOut[12] = fifoOut[14][2][w-1];
              unloadMuxOut[13] = fifoOut[15][2][w-1];
              unloadMuxOut[14] = fifoOut[16][2][w-1];
              unloadMuxOut[15] = fifoOut[17][2][w-1];
              unloadMuxOut[16] = fifoOut[18][2][w-1];
              unloadMuxOut[17] = fifoOut[19][2][w-1];
              unloadMuxOut[18] = fifoOut[20][2][w-1];
              unloadMuxOut[19] = fifoOut[21][2][w-1];
              unloadMuxOut[20] = fifoOut[22][2][w-1];
              unloadMuxOut[21] = fifoOut[23][2][w-1];
              unloadMuxOut[22] = fifoOut[24][2][w-1];
              unloadMuxOut[23] = fifoOut[25][2][w-1];
              unloadMuxOut[24] = fifoOut[0][1][w-1];
              unloadMuxOut[25] = fifoOut[1][1][w-1];
              unloadMuxOut[26] = fifoOut[2][1][w-1];
              unloadMuxOut[27] = fifoOut[3][1][w-1];
              unloadMuxOut[28] = fifoOut[4][1][w-1];
              unloadMuxOut[29] = fifoOut[5][1][w-1];
              unloadMuxOut[30] = fifoOut[6][1][w-1];
              unloadMuxOut[31] = fifoOut[7][1][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[8][1][w-1];
              unloadMuxOut[1] = fifoOut[9][1][w-1];
              unloadMuxOut[2] = fifoOut[10][1][w-1];
              unloadMuxOut[3] = fifoOut[11][1][w-1];
              unloadMuxOut[4] = fifoOut[12][1][w-1];
              unloadMuxOut[5] = fifoOut[13][1][w-1];
              unloadMuxOut[6] = fifoOut[14][1][w-1];
              unloadMuxOut[7] = fifoOut[15][1][w-1];
              unloadMuxOut[8] = fifoOut[16][1][w-1];
              unloadMuxOut[9] = fifoOut[17][1][w-1];
              unloadMuxOut[10] = fifoOut[18][1][w-1];
              unloadMuxOut[11] = fifoOut[19][1][w-1];
              unloadMuxOut[12] = fifoOut[20][1][w-1];
              unloadMuxOut[13] = fifoOut[21][1][w-1];
              unloadMuxOut[14] = fifoOut[22][1][w-1];
              unloadMuxOut[15] = fifoOut[23][1][w-1];
              unloadMuxOut[16] = fifoOut[24][1][w-1];
              unloadMuxOut[17] = fifoOut[25][1][w-1];
              unloadMuxOut[18] = fifoOut[0][0][w-1];
              unloadMuxOut[19] = fifoOut[1][0][w-1];
              unloadMuxOut[20] = fifoOut[2][0][w-1];
              unloadMuxOut[21] = fifoOut[3][0][w-1];
              unloadMuxOut[22] = fifoOut[4][0][w-1];
              unloadMuxOut[23] = fifoOut[5][0][w-1];
              unloadMuxOut[24] = fifoOut[6][0][w-1];
              unloadMuxOut[25] = fifoOut[7][0][w-1];
              unloadMuxOut[26] = fifoOut[26][14][w-1];
              unloadMuxOut[27] = fifoOut[27][14][w-1];
              unloadMuxOut[28] = fifoOut[28][14][w-1];
              unloadMuxOut[29] = fifoOut[29][14][w-1];
              unloadMuxOut[30] = fifoOut[30][14][w-1];
              unloadMuxOut[31] = fifoOut[31][14][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[32][14][w-1];
              unloadMuxOut[1] = fifoOut[33][14][w-1];
              unloadMuxOut[2] = fifoOut[34][14][w-1];
              unloadMuxOut[3] = fifoOut[35][14][w-1];
              unloadMuxOut[4] = fifoOut[36][14][w-1];
              unloadMuxOut[5] = fifoOut[37][14][w-1];
              unloadMuxOut[6] = fifoOut[38][14][w-1];
              unloadMuxOut[7] = fifoOut[39][14][w-1];
              unloadMuxOut[8] = fifoOut[40][14][w-1];
              unloadMuxOut[9] = fifoOut[41][14][w-1];
              unloadMuxOut[10] = fifoOut[42][14][w-1];
              unloadMuxOut[11] = fifoOut[43][14][w-1];
              unloadMuxOut[12] = fifoOut[44][14][w-1];
              unloadMuxOut[13] = fifoOut[45][14][w-1];
              unloadMuxOut[14] = fifoOut[46][14][w-1];
              unloadMuxOut[15] = fifoOut[47][14][w-1];
              unloadMuxOut[16] = fifoOut[48][14][w-1];
              unloadMuxOut[17] = fifoOut[49][14][w-1];
              unloadMuxOut[18] = fifoOut[50][14][w-1];
              unloadMuxOut[19] = fifoOut[51][14][w-1];
              unloadMuxOut[20] = fifoOut[26][13][w-1];
              unloadMuxOut[21] = fifoOut[27][13][w-1];
              unloadMuxOut[22] = fifoOut[28][13][w-1];
              unloadMuxOut[23] = fifoOut[29][13][w-1];
              unloadMuxOut[24] = fifoOut[30][13][w-1];
              unloadMuxOut[25] = fifoOut[31][13][w-1];
              unloadMuxOut[26] = fifoOut[32][13][w-1];
              unloadMuxOut[27] = fifoOut[33][13][w-1];
              unloadMuxOut[28] = fifoOut[34][13][w-1];
              unloadMuxOut[29] = fifoOut[35][13][w-1];
              unloadMuxOut[30] = fifoOut[36][13][w-1];
              unloadMuxOut[31] = fifoOut[37][13][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[38][13][w-1];
              unloadMuxOut[1] = fifoOut[39][13][w-1];
              unloadMuxOut[2] = fifoOut[40][13][w-1];
              unloadMuxOut[3] = fifoOut[41][13][w-1];
              unloadMuxOut[4] = fifoOut[42][13][w-1];
              unloadMuxOut[5] = fifoOut[43][13][w-1];
              unloadMuxOut[6] = fifoOut[44][13][w-1];
              unloadMuxOut[7] = fifoOut[45][13][w-1];
              unloadMuxOut[8] = fifoOut[46][13][w-1];
              unloadMuxOut[9] = fifoOut[47][13][w-1];
              unloadMuxOut[10] = fifoOut[48][13][w-1];
              unloadMuxOut[11] = fifoOut[49][13][w-1];
              unloadMuxOut[12] = fifoOut[50][13][w-1];
              unloadMuxOut[13] = fifoOut[51][13][w-1];
              unloadMuxOut[14] = fifoOut[26][12][w-1];
              unloadMuxOut[15] = fifoOut[27][12][w-1];
              unloadMuxOut[16] = fifoOut[28][12][w-1];
              unloadMuxOut[17] = fifoOut[29][12][w-1];
              unloadMuxOut[18] = fifoOut[30][12][w-1];
              unloadMuxOut[19] = fifoOut[31][12][w-1];
              unloadMuxOut[20] = fifoOut[32][12][w-1];
              unloadMuxOut[21] = fifoOut[33][12][w-1];
              unloadMuxOut[22] = fifoOut[34][12][w-1];
              unloadMuxOut[23] = fifoOut[35][12][w-1];
              unloadMuxOut[24] = fifoOut[36][12][w-1];
              unloadMuxOut[25] = fifoOut[37][12][w-1];
              unloadMuxOut[26] = fifoOut[38][12][w-1];
              unloadMuxOut[27] = fifoOut[39][12][w-1];
              unloadMuxOut[28] = fifoOut[40][12][w-1];
              unloadMuxOut[29] = fifoOut[41][12][w-1];
              unloadMuxOut[30] = fifoOut[42][12][w-1];
              unloadMuxOut[31] = fifoOut[43][12][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[44][12][w-1];
              unloadMuxOut[1] = fifoOut[45][12][w-1];
              unloadMuxOut[2] = fifoOut[46][12][w-1];
              unloadMuxOut[3] = fifoOut[47][12][w-1];
              unloadMuxOut[4] = fifoOut[48][12][w-1];
              unloadMuxOut[5] = fifoOut[49][12][w-1];
              unloadMuxOut[6] = fifoOut[50][12][w-1];
              unloadMuxOut[7] = fifoOut[51][12][w-1];
              unloadMuxOut[8] = fifoOut[26][11][w-1];
              unloadMuxOut[9] = fifoOut[27][11][w-1];
              unloadMuxOut[10] = fifoOut[28][11][w-1];
              unloadMuxOut[11] = fifoOut[29][11][w-1];
              unloadMuxOut[12] = fifoOut[30][11][w-1];
              unloadMuxOut[13] = fifoOut[31][11][w-1];
              unloadMuxOut[14] = fifoOut[32][11][w-1];
              unloadMuxOut[15] = fifoOut[33][11][w-1];
              unloadMuxOut[16] = fifoOut[34][11][w-1];
              unloadMuxOut[17] = fifoOut[35][11][w-1];
              unloadMuxOut[18] = fifoOut[36][11][w-1];
              unloadMuxOut[19] = fifoOut[37][11][w-1];
              unloadMuxOut[20] = fifoOut[38][11][w-1];
              unloadMuxOut[21] = fifoOut[39][11][w-1];
              unloadMuxOut[22] = fifoOut[40][11][w-1];
              unloadMuxOut[23] = fifoOut[41][11][w-1];
              unloadMuxOut[24] = fifoOut[42][11][w-1];
              unloadMuxOut[25] = fifoOut[43][11][w-1];
              unloadMuxOut[26] = fifoOut[44][11][w-1];
              unloadMuxOut[27] = fifoOut[45][11][w-1];
              unloadMuxOut[28] = fifoOut[46][11][w-1];
              unloadMuxOut[29] = fifoOut[47][11][w-1];
              unloadMuxOut[30] = fifoOut[48][11][w-1];
              unloadMuxOut[31] = fifoOut[49][11][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[50][11][w-1];
              unloadMuxOut[1] = fifoOut[51][11][w-1];
              unloadMuxOut[2] = fifoOut[26][10][w-1];
              unloadMuxOut[3] = fifoOut[27][10][w-1];
              unloadMuxOut[4] = fifoOut[28][10][w-1];
              unloadMuxOut[5] = fifoOut[29][10][w-1];
              unloadMuxOut[6] = fifoOut[30][10][w-1];
              unloadMuxOut[7] = fifoOut[31][10][w-1];
              unloadMuxOut[8] = fifoOut[32][10][w-1];
              unloadMuxOut[9] = fifoOut[33][10][w-1];
              unloadMuxOut[10] = fifoOut[34][10][w-1];
              unloadMuxOut[11] = fifoOut[35][10][w-1];
              unloadMuxOut[12] = fifoOut[36][10][w-1];
              unloadMuxOut[13] = fifoOut[37][10][w-1];
              unloadMuxOut[14] = fifoOut[38][10][w-1];
              unloadMuxOut[15] = fifoOut[39][10][w-1];
              unloadMuxOut[16] = fifoOut[40][10][w-1];
              unloadMuxOut[17] = fifoOut[41][10][w-1];
              unloadMuxOut[18] = fifoOut[42][10][w-1];
              unloadMuxOut[19] = fifoOut[43][10][w-1];
              unloadMuxOut[20] = fifoOut[44][10][w-1];
              unloadMuxOut[21] = fifoOut[45][10][w-1];
              unloadMuxOut[22] = fifoOut[46][10][w-1];
              unloadMuxOut[23] = fifoOut[47][10][w-1];
              unloadMuxOut[24] = fifoOut[48][10][w-1];
              unloadMuxOut[25] = fifoOut[49][10][w-1];
              unloadMuxOut[26] = fifoOut[50][10][w-1];
              unloadMuxOut[27] = fifoOut[51][10][w-1];
              unloadMuxOut[28] = fifoOut[26][9][w-1];
              unloadMuxOut[29] = fifoOut[27][9][w-1];
              unloadMuxOut[30] = fifoOut[28][9][w-1];
              unloadMuxOut[31] = fifoOut[29][9][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[30][9][w-1];
              unloadMuxOut[1] = fifoOut[31][9][w-1];
              unloadMuxOut[2] = fifoOut[32][9][w-1];
              unloadMuxOut[3] = fifoOut[33][9][w-1];
              unloadMuxOut[4] = fifoOut[34][9][w-1];
              unloadMuxOut[5] = fifoOut[0][14][w-1];
              unloadMuxOut[6] = fifoOut[1][14][w-1];
              unloadMuxOut[7] = fifoOut[2][14][w-1];
              unloadMuxOut[8] = fifoOut[3][14][w-1];
              unloadMuxOut[9] = fifoOut[4][14][w-1];
              unloadMuxOut[10] = fifoOut[5][14][w-1];
              unloadMuxOut[11] = fifoOut[6][14][w-1];
              unloadMuxOut[12] = fifoOut[7][14][w-1];
              unloadMuxOut[13] = fifoOut[8][14][w-1];
              unloadMuxOut[14] = fifoOut[9][14][w-1];
              unloadMuxOut[15] = fifoOut[10][14][w-1];
              unloadMuxOut[16] = fifoOut[11][14][w-1];
              unloadMuxOut[17] = fifoOut[12][14][w-1];
              unloadMuxOut[18] = fifoOut[13][14][w-1];
              unloadMuxOut[19] = fifoOut[14][14][w-1];
              unloadMuxOut[20] = fifoOut[15][14][w-1];
              unloadMuxOut[21] = fifoOut[16][14][w-1];
              unloadMuxOut[22] = fifoOut[17][14][w-1];
              unloadMuxOut[23] = fifoOut[18][14][w-1];
              unloadMuxOut[24] = fifoOut[19][14][w-1];
              unloadMuxOut[25] = fifoOut[20][14][w-1];
              unloadMuxOut[26] = fifoOut[21][14][w-1];
              unloadMuxOut[27] = fifoOut[22][14][w-1];
              unloadMuxOut[28] = fifoOut[23][14][w-1];
              unloadMuxOut[29] = fifoOut[24][14][w-1];
              unloadMuxOut[30] = fifoOut[25][14][w-1];
              unloadMuxOut[31] = fifoOut[0][13][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[1][13][w-1];
              unloadMuxOut[1] = fifoOut[2][13][w-1];
              unloadMuxOut[2] = fifoOut[3][13][w-1];
              unloadMuxOut[3] = fifoOut[4][13][w-1];
              unloadMuxOut[4] = fifoOut[5][13][w-1];
              unloadMuxOut[5] = fifoOut[6][13][w-1];
              unloadMuxOut[6] = fifoOut[7][13][w-1];
              unloadMuxOut[7] = fifoOut[8][13][w-1];
              unloadMuxOut[8] = fifoOut[9][13][w-1];
              unloadMuxOut[9] = fifoOut[10][13][w-1];
              unloadMuxOut[10] = fifoOut[11][13][w-1];
              unloadMuxOut[11] = fifoOut[12][13][w-1];
              unloadMuxOut[12] = fifoOut[13][13][w-1];
              unloadMuxOut[13] = fifoOut[14][13][w-1];
              unloadMuxOut[14] = fifoOut[15][13][w-1];
              unloadMuxOut[15] = fifoOut[16][13][w-1];
              unloadMuxOut[16] = fifoOut[17][13][w-1];
              unloadMuxOut[17] = fifoOut[18][13][w-1];
              unloadMuxOut[18] = fifoOut[19][13][w-1];
              unloadMuxOut[19] = fifoOut[20][13][w-1];
              unloadMuxOut[20] = fifoOut[21][13][w-1];
              unloadMuxOut[21] = fifoOut[22][13][w-1];
              unloadMuxOut[22] = fifoOut[23][13][w-1];
              unloadMuxOut[23] = fifoOut[24][13][w-1];
              unloadMuxOut[24] = fifoOut[25][13][w-1];
              unloadMuxOut[25] = fifoOut[0][12][w-1];
              unloadMuxOut[26] = fifoOut[1][12][w-1];
              unloadMuxOut[27] = fifoOut[2][12][w-1];
              unloadMuxOut[28] = fifoOut[3][12][w-1];
              unloadMuxOut[29] = fifoOut[4][12][w-1];
              unloadMuxOut[30] = fifoOut[5][12][w-1];
              unloadMuxOut[31] = fifoOut[6][12][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[7][12][w-1];
              unloadMuxOut[1] = fifoOut[8][12][w-1];
              unloadMuxOut[2] = fifoOut[9][12][w-1];
              unloadMuxOut[3] = fifoOut[10][12][w-1];
              unloadMuxOut[4] = fifoOut[11][12][w-1];
              unloadMuxOut[5] = fifoOut[12][12][w-1];
              unloadMuxOut[6] = fifoOut[13][12][w-1];
              unloadMuxOut[7] = fifoOut[14][12][w-1];
              unloadMuxOut[8] = fifoOut[15][12][w-1];
              unloadMuxOut[9] = fifoOut[16][12][w-1];
              unloadMuxOut[10] = fifoOut[17][12][w-1];
              unloadMuxOut[11] = fifoOut[18][12][w-1];
              unloadMuxOut[12] = fifoOut[19][12][w-1];
              unloadMuxOut[13] = fifoOut[20][12][w-1];
              unloadMuxOut[14] = fifoOut[21][12][w-1];
              unloadMuxOut[15] = fifoOut[22][12][w-1];
              unloadMuxOut[16] = fifoOut[23][12][w-1];
              unloadMuxOut[17] = fifoOut[24][12][w-1];
              unloadMuxOut[18] = fifoOut[25][12][w-1];
              unloadMuxOut[19] = fifoOut[0][11][w-1];
              unloadMuxOut[20] = fifoOut[1][11][w-1];
              unloadMuxOut[21] = fifoOut[2][11][w-1];
              unloadMuxOut[22] = fifoOut[3][11][w-1];
              unloadMuxOut[23] = fifoOut[4][11][w-1];
              unloadMuxOut[24] = fifoOut[5][11][w-1];
              unloadMuxOut[25] = fifoOut[6][11][w-1];
              unloadMuxOut[26] = fifoOut[7][11][w-1];
              unloadMuxOut[27] = fifoOut[8][11][w-1];
              unloadMuxOut[28] = fifoOut[9][11][w-1];
              unloadMuxOut[29] = fifoOut[10][11][w-1];
              unloadMuxOut[30] = fifoOut[11][11][w-1];
              unloadMuxOut[31] = fifoOut[12][11][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[13][11][w-1];
              unloadMuxOut[1] = fifoOut[14][11][w-1];
              unloadMuxOut[2] = fifoOut[15][11][w-1];
              unloadMuxOut[3] = fifoOut[16][11][w-1];
              unloadMuxOut[4] = fifoOut[17][11][w-1];
              unloadMuxOut[5] = fifoOut[18][11][w-1];
              unloadMuxOut[6] = fifoOut[19][11][w-1];
              unloadMuxOut[7] = fifoOut[20][11][w-1];
              unloadMuxOut[8] = fifoOut[21][11][w-1];
              unloadMuxOut[9] = fifoOut[22][11][w-1];
              unloadMuxOut[10] = fifoOut[23][11][w-1];
              unloadMuxOut[11] = fifoOut[24][11][w-1];
              unloadMuxOut[12] = fifoOut[25][11][w-1];
              unloadMuxOut[13] = fifoOut[0][10][w-1];
              unloadMuxOut[14] = fifoOut[1][10][w-1];
              unloadMuxOut[15] = fifoOut[2][10][w-1];
              unloadMuxOut[16] = fifoOut[3][10][w-1];
              unloadMuxOut[17] = fifoOut[4][10][w-1];
              unloadMuxOut[18] = fifoOut[5][10][w-1];
              unloadMuxOut[19] = fifoOut[6][10][w-1];
              unloadMuxOut[20] = fifoOut[7][10][w-1];
              unloadMuxOut[21] = fifoOut[8][10][w-1];
              unloadMuxOut[22] = fifoOut[9][10][w-1];
              unloadMuxOut[23] = fifoOut[10][10][w-1];
              unloadMuxOut[24] = fifoOut[11][10][w-1];
              unloadMuxOut[25] = fifoOut[12][10][w-1];
              unloadMuxOut[26] = fifoOut[13][10][w-1];
              unloadMuxOut[27] = fifoOut[14][10][w-1];
              unloadMuxOut[28] = fifoOut[15][10][w-1];
              unloadMuxOut[29] = fifoOut[16][10][w-1];
              unloadMuxOut[30] = fifoOut[17][10][w-1];
              unloadMuxOut[31] = fifoOut[18][10][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[19][10][w-1];
              unloadMuxOut[1] = fifoOut[20][10][w-1];
              unloadMuxOut[2] = fifoOut[21][10][w-1];
              unloadMuxOut[3] = fifoOut[22][10][w-1];
              unloadMuxOut[4] = fifoOut[23][10][w-1];
              unloadMuxOut[5] = fifoOut[24][10][w-1];
              unloadMuxOut[6] = fifoOut[25][10][w-1];
              unloadMuxOut[7] = fifoOut[0][9][w-1];
              unloadMuxOut[8] = fifoOut[1][9][w-1];
              unloadMuxOut[9] = fifoOut[2][9][w-1];
              unloadMuxOut[10] = fifoOut[3][9][w-1];
              unloadMuxOut[11] = fifoOut[4][9][w-1];
              unloadMuxOut[12] = fifoOut[5][9][w-1];
              unloadMuxOut[13] = fifoOut[6][9][w-1];
              unloadMuxOut[14] = fifoOut[7][9][w-1];
              unloadMuxOut[15] = fifoOut[8][9][w-1];
              unloadMuxOut[16] = fifoOut[9][9][w-1];
              unloadMuxOut[17] = fifoOut[10][9][w-1];
              unloadMuxOut[18] = fifoOut[11][9][w-1];
              unloadMuxOut[19] = fifoOut[12][9][w-1];
              unloadMuxOut[20] = fifoOut[13][9][w-1];
              unloadMuxOut[21] = fifoOut[14][9][w-1];
              unloadMuxOut[22] = fifoOut[15][9][w-1];
              unloadMuxOut[23] = fifoOut[16][9][w-1];
              unloadMuxOut[24] = fifoOut[17][9][w-1];
              unloadMuxOut[25] = fifoOut[18][9][w-1];
              unloadMuxOut[26] = fifoOut[19][9][w-1];
              unloadMuxOut[27] = fifoOut[20][9][w-1];
              unloadMuxOut[28] = fifoOut[21][9][w-1];
              unloadMuxOut[29] = fifoOut[22][9][w-1];
              unloadMuxOut[30] = fifoOut[23][9][w-1];
              unloadMuxOut[31] = fifoOut[24][9][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[25][9][w-1];
              unloadMuxOut[1] = fifoOut[0][8][w-1];
              unloadMuxOut[2] = fifoOut[1][8][w-1];
              unloadMuxOut[3] = fifoOut[2][8][w-1];
              unloadMuxOut[4] = fifoOut[3][8][w-1];
              unloadMuxOut[5] = fifoOut[4][8][w-1];
              unloadMuxOut[6] = fifoOut[5][8][w-1];
              unloadMuxOut[7] = fifoOut[6][8][w-1];
              unloadMuxOut[8] = fifoOut[7][8][w-1];
              unloadMuxOut[9] = fifoOut[8][8][w-1];
              unloadMuxOut[10] = fifoOut[9][8][w-1];
              unloadMuxOut[11] = fifoOut[10][8][w-1];
              unloadMuxOut[12] = fifoOut[11][8][w-1];
              unloadMuxOut[13] = fifoOut[12][8][w-1];
              unloadMuxOut[14] = fifoOut[13][8][w-1];
              unloadMuxOut[15] = fifoOut[14][8][w-1];
              unloadMuxOut[16] = fifoOut[15][8][w-1];
              unloadMuxOut[17] = fifoOut[16][8][w-1];
              unloadMuxOut[18] = fifoOut[17][8][w-1];
              unloadMuxOut[19] = fifoOut[18][8][w-1];
              unloadMuxOut[20] = fifoOut[19][8][w-1];
              unloadMuxOut[21] = fifoOut[20][8][w-1];
              unloadMuxOut[22] = fifoOut[21][8][w-1];
              unloadMuxOut[23] = fifoOut[22][8][w-1];
              unloadMuxOut[24] = fifoOut[23][8][w-1];
              unloadMuxOut[25] = fifoOut[24][8][w-1];
              unloadMuxOut[26] = fifoOut[25][8][w-1];
              unloadMuxOut[27] = fifoOut[0][7][w-1];
              unloadMuxOut[28] = fifoOut[1][7][w-1];
              unloadMuxOut[29] = fifoOut[2][7][w-1];
              unloadMuxOut[30] = fifoOut[3][7][w-1];
              unloadMuxOut[31] = fifoOut[4][7][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[5][7][w-1];
              unloadMuxOut[1] = fifoOut[6][7][w-1];
              unloadMuxOut[2] = fifoOut[7][7][w-1];
              unloadMuxOut[3] = fifoOut[8][7][w-1];
              unloadMuxOut[4] = fifoOut[9][7][w-1];
              unloadMuxOut[5] = fifoOut[10][7][w-1];
              unloadMuxOut[6] = fifoOut[11][7][w-1];
              unloadMuxOut[7] = fifoOut[12][7][w-1];
              unloadMuxOut[8] = fifoOut[13][7][w-1];
              unloadMuxOut[9] = fifoOut[14][7][w-1];
              unloadMuxOut[10] = fifoOut[15][7][w-1];
              unloadMuxOut[11] = fifoOut[16][7][w-1];
              unloadMuxOut[12] = fifoOut[17][7][w-1];
              unloadMuxOut[13] = fifoOut[18][7][w-1];
              unloadMuxOut[14] = fifoOut[19][7][w-1];
              unloadMuxOut[15] = fifoOut[20][7][w-1];
              unloadMuxOut[16] = fifoOut[21][7][w-1];
              unloadMuxOut[17] = fifoOut[22][7][w-1];
              unloadMuxOut[18] = fifoOut[23][7][w-1];
              unloadMuxOut[19] = fifoOut[24][7][w-1];
              unloadMuxOut[20] = fifoOut[25][7][w-1];
              unloadMuxOut[21] = fifoOut[0][6][w-1];
              unloadMuxOut[22] = fifoOut[1][6][w-1];
              unloadMuxOut[23] = fifoOut[2][6][w-1];
              unloadMuxOut[24] = fifoOut[3][6][w-1];
              unloadMuxOut[25] = fifoOut[4][6][w-1];
              unloadMuxOut[26] = fifoOut[5][6][w-1];
              unloadMuxOut[27] = fifoOut[6][6][w-1];
              unloadMuxOut[28] = fifoOut[7][6][w-1];
              unloadMuxOut[29] = fifoOut[8][6][w-1];
              unloadMuxOut[30] = fifoOut[9][6][w-1];
              unloadMuxOut[31] = fifoOut[10][6][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[11][6][w-1];
              unloadMuxOut[1] = fifoOut[12][6][w-1];
              unloadMuxOut[2] = fifoOut[13][6][w-1];
              unloadMuxOut[3] = fifoOut[14][6][w-1];
              unloadMuxOut[4] = fifoOut[15][6][w-1];
              unloadMuxOut[5] = fifoOut[16][6][w-1];
              unloadMuxOut[6] = fifoOut[17][6][w-1];
              unloadMuxOut[7] = fifoOut[18][6][w-1];
              unloadMuxOut[8] = fifoOut[19][6][w-1];
              unloadMuxOut[9] = fifoOut[20][6][w-1];
              unloadMuxOut[10] = fifoOut[21][6][w-1];
              unloadMuxOut[11] = fifoOut[22][6][w-1];
              unloadMuxOut[12] = fifoOut[23][6][w-1];
              unloadMuxOut[13] = fifoOut[24][6][w-1];
              unloadMuxOut[14] = fifoOut[25][6][w-1];
              unloadMuxOut[15] = fifoOut[0][5][w-1];
              unloadMuxOut[16] = fifoOut[1][5][w-1];
              unloadMuxOut[17] = fifoOut[2][5][w-1];
              unloadMuxOut[18] = fifoOut[3][5][w-1];
              unloadMuxOut[19] = fifoOut[4][5][w-1];
              unloadMuxOut[20] = fifoOut[5][5][w-1];
              unloadMuxOut[21] = fifoOut[6][5][w-1];
              unloadMuxOut[22] = fifoOut[7][5][w-1];
              unloadMuxOut[23] = fifoOut[8][5][w-1];
              unloadMuxOut[24] = fifoOut[9][5][w-1];
              unloadMuxOut[25] = fifoOut[10][5][w-1];
              unloadMuxOut[26] = fifoOut[11][5][w-1];
              unloadMuxOut[27] = fifoOut[12][5][w-1];
              unloadMuxOut[28] = fifoOut[13][5][w-1];
              unloadMuxOut[29] = fifoOut[14][5][w-1];
              unloadMuxOut[30] = fifoOut[15][5][w-1];
              unloadMuxOut[31] = fifoOut[16][5][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[17][5][w-1];
              unloadMuxOut[1] = fifoOut[18][5][w-1];
              unloadMuxOut[2] = fifoOut[19][5][w-1];
              unloadMuxOut[3] = fifoOut[20][5][w-1];
              unloadMuxOut[4] = fifoOut[21][5][w-1];
              unloadMuxOut[5] = fifoOut[22][5][w-1];
              unloadMuxOut[6] = fifoOut[23][5][w-1];
              unloadMuxOut[7] = fifoOut[24][5][w-1];
              unloadMuxOut[8] = fifoOut[25][5][w-1];
              unloadMuxOut[9] = fifoOut[0][4][w-1];
              unloadMuxOut[10] = fifoOut[1][4][w-1];
              unloadMuxOut[11] = fifoOut[2][4][w-1];
              unloadMuxOut[12] = fifoOut[3][4][w-1];
              unloadMuxOut[13] = fifoOut[4][4][w-1];
              unloadMuxOut[14] = fifoOut[5][4][w-1];
              unloadMuxOut[15] = fifoOut[6][4][w-1];
              unloadMuxOut[16] = fifoOut[7][4][w-1];
              unloadMuxOut[17] = fifoOut[8][4][w-1];
              unloadMuxOut[18] = fifoOut[9][4][w-1];
              unloadMuxOut[19] = fifoOut[10][4][w-1];
              unloadMuxOut[20] = fifoOut[11][4][w-1];
              unloadMuxOut[21] = fifoOut[12][4][w-1];
              unloadMuxOut[22] = fifoOut[13][4][w-1];
              unloadMuxOut[23] = fifoOut[14][4][w-1];
              unloadMuxOut[24] = fifoOut[15][4][w-1];
              unloadMuxOut[25] = fifoOut[16][4][w-1];
              unloadMuxOut[26] = fifoOut[17][4][w-1];
              unloadMuxOut[27] = fifoOut[18][4][w-1];
              unloadMuxOut[28] = fifoOut[19][4][w-1];
              unloadMuxOut[29] = fifoOut[20][4][w-1];
              unloadMuxOut[30] = fifoOut[21][4][w-1];
              unloadMuxOut[31] = 1'b0;
       end
       16: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0;
             end
       end
    endcase
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[22][4];
              muxOutConnector[1] = fifoOut[23][4];
              muxOutConnector[2] = fifoOut[24][4];
              muxOutConnector[3] = fifoOut[25][4];
              muxOutConnector[4] = fifoOut[0][3];
              muxOutConnector[5] = fifoOut[1][3];
              muxOutConnector[6] = fifoOut[2][3];
              muxOutConnector[7] = fifoOut[3][3];
              muxOutConnector[8] = fifoOut[4][3];
              muxOutConnector[9] = fifoOut[5][3];
              muxOutConnector[10] = fifoOut[6][3];
              muxOutConnector[11] = fifoOut[7][3];
              muxOutConnector[12] = fifoOut[8][3];
              muxOutConnector[13] = fifoOut[9][3];
              muxOutConnector[14] = fifoOut[10][3];
              muxOutConnector[15] = fifoOut[11][3];
              muxOutConnector[16] = fifoOut[12][3];
              muxOutConnector[17] = fifoOut[13][3];
              muxOutConnector[18] = fifoOut[14][3];
              muxOutConnector[19] = fifoOut[15][3];
              muxOutConnector[20] = fifoOut[16][3];
              muxOutConnector[21] = fifoOut[17][3];
              muxOutConnector[22] = fifoOut[18][3];
              muxOutConnector[23] = fifoOut[19][3];
              muxOutConnector[24] = fifoOut[20][3];
              muxOutConnector[25] = fifoOut[21][3];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[35][11];
              muxOutConnector[28] = fifoOut[36][11];
              muxOutConnector[29] = fifoOut[37][11];
              muxOutConnector[30] = fifoOut[38][11];
              muxOutConnector[31] = fifoOut[39][11];
              muxOutConnector[32] = fifoOut[40][11];
              muxOutConnector[33] = fifoOut[41][11];
              muxOutConnector[34] = fifoOut[42][11];
              muxOutConnector[35] = fifoOut[43][11];
              muxOutConnector[36] = fifoOut[44][11];
              muxOutConnector[37] = fifoOut[45][11];
              muxOutConnector[38] = fifoOut[46][11];
              muxOutConnector[39] = fifoOut[47][11];
              muxOutConnector[40] = fifoOut[48][11];
              muxOutConnector[41] = fifoOut[49][11];
              muxOutConnector[42] = fifoOut[50][11];
              muxOutConnector[43] = fifoOut[51][11];
              muxOutConnector[44] = fifoOut[26][10];
              muxOutConnector[45] = fifoOut[27][10];
              muxOutConnector[46] = fifoOut[28][10];
              muxOutConnector[47] = fifoOut[29][10];
              muxOutConnector[48] = fifoOut[30][10];
              muxOutConnector[49] = fifoOut[31][10];
              muxOutConnector[50] = fifoOut[32][10];
              muxOutConnector[51] = fifoOut[33][10];
       end
       1: begin
              muxOutConnector[0] = fifoOut[22][4];
              muxOutConnector[1] = fifoOut[23][4];
              muxOutConnector[2] = fifoOut[24][4];
              muxOutConnector[3] = fifoOut[25][4];
              muxOutConnector[4] = fifoOut[0][3];
              muxOutConnector[5] = fifoOut[1][3];
              muxOutConnector[6] = fifoOut[2][3];
              muxOutConnector[7] = fifoOut[3][3];
              muxOutConnector[8] = fifoOut[4][3];
              muxOutConnector[9] = fifoOut[5][3];
              muxOutConnector[10] = fifoOut[6][3];
              muxOutConnector[11] = fifoOut[7][3];
              muxOutConnector[12] = fifoOut[8][3];
              muxOutConnector[13] = fifoOut[9][3];
              muxOutConnector[14] = fifoOut[10][3];
              muxOutConnector[15] = fifoOut[11][3];
              muxOutConnector[16] = fifoOut[12][3];
              muxOutConnector[17] = fifoOut[13][3];
              muxOutConnector[18] = fifoOut[14][3];
              muxOutConnector[19] = fifoOut[15][3];
              muxOutConnector[20] = fifoOut[16][3];
              muxOutConnector[21] = fifoOut[17][3];
              muxOutConnector[22] = fifoOut[18][3];
              muxOutConnector[23] = fifoOut[19][3];
              muxOutConnector[24] = fifoOut[20][3];
              muxOutConnector[25] = fifoOut[21][3];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[35][11];
              muxOutConnector[28] = fifoOut[36][11];
              muxOutConnector[29] = fifoOut[37][11];
              muxOutConnector[30] = fifoOut[38][11];
              muxOutConnector[31] = fifoOut[39][11];
              muxOutConnector[32] = fifoOut[40][11];
              muxOutConnector[33] = fifoOut[41][11];
              muxOutConnector[34] = fifoOut[42][11];
              muxOutConnector[35] = fifoOut[43][11];
              muxOutConnector[36] = fifoOut[44][11];
              muxOutConnector[37] = fifoOut[45][11];
              muxOutConnector[38] = fifoOut[46][11];
              muxOutConnector[39] = fifoOut[47][11];
              muxOutConnector[40] = fifoOut[48][11];
              muxOutConnector[41] = fifoOut[49][11];
              muxOutConnector[42] = fifoOut[50][11];
              muxOutConnector[43] = fifoOut[51][11];
              muxOutConnector[44] = fifoOut[26][10];
              muxOutConnector[45] = fifoOut[27][10];
              muxOutConnector[46] = fifoOut[28][10];
              muxOutConnector[47] = fifoOut[29][10];
              muxOutConnector[48] = fifoOut[30][10];
              muxOutConnector[49] = fifoOut[31][10];
              muxOutConnector[50] = fifoOut[32][10];
              muxOutConnector[51] = fifoOut[33][10];
       end
       2: begin
              muxOutConnector[0] = fifoOut[22][4];
              muxOutConnector[1] = fifoOut[23][4];
              muxOutConnector[2] = fifoOut[24][4];
              muxOutConnector[3] = fifoOut[25][4];
              muxOutConnector[4] = fifoOut[0][3];
              muxOutConnector[5] = fifoOut[1][3];
              muxOutConnector[6] = fifoOut[2][3];
              muxOutConnector[7] = fifoOut[3][3];
              muxOutConnector[8] = fifoOut[4][3];
              muxOutConnector[9] = fifoOut[5][3];
              muxOutConnector[10] = fifoOut[6][3];
              muxOutConnector[11] = fifoOut[7][3];
              muxOutConnector[12] = fifoOut[8][3];
              muxOutConnector[13] = fifoOut[9][3];
              muxOutConnector[14] = fifoOut[10][3];
              muxOutConnector[15] = fifoOut[11][3];
              muxOutConnector[16] = fifoOut[12][3];
              muxOutConnector[17] = fifoOut[13][3];
              muxOutConnector[18] = fifoOut[14][3];
              muxOutConnector[19] = fifoOut[15][3];
              muxOutConnector[20] = fifoOut[16][3];
              muxOutConnector[21] = fifoOut[17][3];
              muxOutConnector[22] = fifoOut[18][3];
              muxOutConnector[23] = fifoOut[19][3];
              muxOutConnector[24] = fifoOut[20][3];
              muxOutConnector[25] = fifoOut[21][3];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[35][11];
              muxOutConnector[28] = fifoOut[36][11];
              muxOutConnector[29] = fifoOut[37][11];
              muxOutConnector[30] = fifoOut[38][11];
              muxOutConnector[31] = fifoOut[39][11];
              muxOutConnector[32] = fifoOut[40][11];
              muxOutConnector[33] = fifoOut[41][11];
              muxOutConnector[34] = fifoOut[42][11];
              muxOutConnector[35] = fifoOut[43][11];
              muxOutConnector[36] = fifoOut[44][11];
              muxOutConnector[37] = fifoOut[45][11];
              muxOutConnector[38] = fifoOut[46][11];
              muxOutConnector[39] = fifoOut[47][11];
              muxOutConnector[40] = fifoOut[48][11];
              muxOutConnector[41] = fifoOut[49][11];
              muxOutConnector[42] = fifoOut[50][11];
              muxOutConnector[43] = fifoOut[51][11];
              muxOutConnector[44] = fifoOut[26][10];
              muxOutConnector[45] = fifoOut[27][10];
              muxOutConnector[46] = fifoOut[28][10];
              muxOutConnector[47] = fifoOut[29][10];
              muxOutConnector[48] = fifoOut[30][10];
              muxOutConnector[49] = fifoOut[31][10];
              muxOutConnector[50] = fifoOut[32][10];
              muxOutConnector[51] = fifoOut[33][10];
       end
       3: begin
              muxOutConnector[0] = fifoOut[22][4];
              muxOutConnector[1] = fifoOut[23][4];
              muxOutConnector[2] = fifoOut[24][4];
              muxOutConnector[3] = fifoOut[25][4];
              muxOutConnector[4] = fifoOut[0][3];
              muxOutConnector[5] = fifoOut[1][3];
              muxOutConnector[6] = fifoOut[2][3];
              muxOutConnector[7] = fifoOut[3][3];
              muxOutConnector[8] = fifoOut[4][3];
              muxOutConnector[9] = fifoOut[5][3];
              muxOutConnector[10] = fifoOut[6][3];
              muxOutConnector[11] = fifoOut[7][3];
              muxOutConnector[12] = fifoOut[8][3];
              muxOutConnector[13] = fifoOut[9][3];
              muxOutConnector[14] = fifoOut[10][3];
              muxOutConnector[15] = fifoOut[11][3];
              muxOutConnector[16] = fifoOut[12][3];
              muxOutConnector[17] = fifoOut[13][3];
              muxOutConnector[18] = fifoOut[14][3];
              muxOutConnector[19] = fifoOut[15][3];
              muxOutConnector[20] = fifoOut[16][3];
              muxOutConnector[21] = fifoOut[35][2];
              muxOutConnector[22] = fifoOut[36][2];
              muxOutConnector[23] = fifoOut[37][2];
              muxOutConnector[24] = fifoOut[38][2];
              muxOutConnector[25] = fifoOut[39][2];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[35][11];
              muxOutConnector[28] = fifoOut[36][11];
              muxOutConnector[29] = fifoOut[37][11];
              muxOutConnector[30] = fifoOut[38][11];
              muxOutConnector[31] = fifoOut[39][11];
              muxOutConnector[32] = fifoOut[40][11];
              muxOutConnector[33] = fifoOut[41][11];
              muxOutConnector[34] = fifoOut[42][11];
              muxOutConnector[35] = fifoOut[43][11];
              muxOutConnector[36] = fifoOut[44][11];
              muxOutConnector[37] = fifoOut[45][11];
              muxOutConnector[38] = fifoOut[46][11];
              muxOutConnector[39] = fifoOut[47][11];
              muxOutConnector[40] = fifoOut[48][11];
              muxOutConnector[41] = fifoOut[49][11];
              muxOutConnector[42] = fifoOut[50][11];
              muxOutConnector[43] = fifoOut[51][11];
              muxOutConnector[44] = fifoOut[26][10];
              muxOutConnector[45] = fifoOut[27][10];
              muxOutConnector[46] = fifoOut[28][10];
              muxOutConnector[47] = fifoOut[29][10];
              muxOutConnector[48] = fifoOut[30][10];
              muxOutConnector[49] = fifoOut[31][10];
              muxOutConnector[50] = fifoOut[32][10];
              muxOutConnector[51] = fifoOut[33][10];
       end
       4: begin
              muxOutConnector[0] = fifoOut[40][3];
              muxOutConnector[1] = fifoOut[41][3];
              muxOutConnector[2] = fifoOut[42][3];
              muxOutConnector[3] = fifoOut[43][3];
              muxOutConnector[4] = fifoOut[44][3];
              muxOutConnector[5] = fifoOut[45][3];
              muxOutConnector[6] = fifoOut[46][3];
              muxOutConnector[7] = fifoOut[47][3];
              muxOutConnector[8] = fifoOut[48][3];
              muxOutConnector[9] = fifoOut[49][3];
              muxOutConnector[10] = fifoOut[50][3];
              muxOutConnector[11] = fifoOut[51][3];
              muxOutConnector[12] = fifoOut[26][2];
              muxOutConnector[13] = fifoOut[27][2];
              muxOutConnector[14] = fifoOut[28][2];
              muxOutConnector[15] = fifoOut[29][2];
              muxOutConnector[16] = fifoOut[30][2];
              muxOutConnector[17] = fifoOut[31][2];
              muxOutConnector[18] = fifoOut[32][2];
              muxOutConnector[19] = fifoOut[33][2];
              muxOutConnector[20] = fifoOut[34][2];
              muxOutConnector[21] = fifoOut[35][2];
              muxOutConnector[22] = fifoOut[36][2];
              muxOutConnector[23] = fifoOut[37][2];
              muxOutConnector[24] = fifoOut[38][2];
              muxOutConnector[25] = fifoOut[39][2];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[35][11];
              muxOutConnector[28] = fifoOut[36][11];
              muxOutConnector[29] = fifoOut[37][11];
              muxOutConnector[30] = fifoOut[38][11];
              muxOutConnector[31] = fifoOut[39][11];
              muxOutConnector[32] = fifoOut[40][11];
              muxOutConnector[33] = fifoOut[41][11];
              muxOutConnector[34] = fifoOut[42][11];
              muxOutConnector[35] = fifoOut[43][11];
              muxOutConnector[36] = fifoOut[44][11];
              muxOutConnector[37] = fifoOut[45][11];
              muxOutConnector[38] = fifoOut[46][11];
              muxOutConnector[39] = fifoOut[47][11];
              muxOutConnector[40] = fifoOut[48][11];
              muxOutConnector[41] = fifoOut[49][11];
              muxOutConnector[42] = fifoOut[50][11];
              muxOutConnector[43] = fifoOut[51][11];
              muxOutConnector[44] = fifoOut[26][10];
              muxOutConnector[45] = fifoOut[27][10];
              muxOutConnector[46] = fifoOut[28][10];
              muxOutConnector[47] = fifoOut[29][10];
              muxOutConnector[48] = fifoOut[30][10];
              muxOutConnector[49] = fifoOut[31][10];
              muxOutConnector[50] = fifoOut[32][10];
              muxOutConnector[51] = fifoOut[33][10];
       end
       5: begin
              muxOutConnector[0] = fifoOut[40][3];
              muxOutConnector[1] = fifoOut[41][3];
              muxOutConnector[2] = fifoOut[42][3];
              muxOutConnector[3] = fifoOut[43][3];
              muxOutConnector[4] = fifoOut[44][3];
              muxOutConnector[5] = fifoOut[45][3];
              muxOutConnector[6] = fifoOut[46][3];
              muxOutConnector[7] = fifoOut[47][3];
              muxOutConnector[8] = fifoOut[48][3];
              muxOutConnector[9] = fifoOut[49][3];
              muxOutConnector[10] = fifoOut[50][3];
              muxOutConnector[11] = fifoOut[51][3];
              muxOutConnector[12] = fifoOut[26][2];
              muxOutConnector[13] = fifoOut[27][2];
              muxOutConnector[14] = fifoOut[28][2];
              muxOutConnector[15] = fifoOut[29][2];
              muxOutConnector[16] = fifoOut[30][2];
              muxOutConnector[17] = fifoOut[31][2];
              muxOutConnector[18] = fifoOut[32][2];
              muxOutConnector[19] = fifoOut[33][2];
              muxOutConnector[20] = fifoOut[34][2];
              muxOutConnector[21] = fifoOut[35][2];
              muxOutConnector[22] = fifoOut[36][2];
              muxOutConnector[23] = fifoOut[37][2];
              muxOutConnector[24] = fifoOut[38][2];
              muxOutConnector[25] = fifoOut[39][2];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[35][11];
              muxOutConnector[28] = fifoOut[36][11];
              muxOutConnector[29] = fifoOut[37][11];
              muxOutConnector[30] = fifoOut[38][11];
              muxOutConnector[31] = fifoOut[39][11];
              muxOutConnector[32] = fifoOut[40][11];
              muxOutConnector[33] = fifoOut[41][11];
              muxOutConnector[34] = fifoOut[42][11];
              muxOutConnector[35] = fifoOut[43][11];
              muxOutConnector[36] = fifoOut[44][11];
              muxOutConnector[37] = fifoOut[45][11];
              muxOutConnector[38] = fifoOut[46][11];
              muxOutConnector[39] = fifoOut[47][11];
              muxOutConnector[40] = fifoOut[48][11];
              muxOutConnector[41] = fifoOut[49][11];
              muxOutConnector[42] = fifoOut[50][11];
              muxOutConnector[43] = fifoOut[51][11];
              muxOutConnector[44] = fifoOut[26][10];
              muxOutConnector[45] = fifoOut[27][10];
              muxOutConnector[46] = fifoOut[28][10];
              muxOutConnector[47] = fifoOut[29][10];
              muxOutConnector[48] = fifoOut[30][10];
              muxOutConnector[49] = fifoOut[31][10];
              muxOutConnector[50] = fifoOut[32][10];
              muxOutConnector[51] = fifoOut[33][10];
       end
       6: begin
              muxOutConnector[0] = fifoOut[40][3];
              muxOutConnector[1] = fifoOut[41][3];
              muxOutConnector[2] = fifoOut[42][3];
              muxOutConnector[3] = fifoOut[43][3];
              muxOutConnector[4] = fifoOut[44][3];
              muxOutConnector[5] = fifoOut[45][3];
              muxOutConnector[6] = fifoOut[46][3];
              muxOutConnector[7] = fifoOut[47][3];
              muxOutConnector[8] = fifoOut[48][3];
              muxOutConnector[9] = fifoOut[49][3];
              muxOutConnector[10] = fifoOut[50][3];
              muxOutConnector[11] = fifoOut[51][3];
              muxOutConnector[12] = fifoOut[26][2];
              muxOutConnector[13] = fifoOut[27][2];
              muxOutConnector[14] = fifoOut[28][2];
              muxOutConnector[15] = fifoOut[29][2];
              muxOutConnector[16] = fifoOut[30][2];
              muxOutConnector[17] = fifoOut[31][2];
              muxOutConnector[18] = fifoOut[32][2];
              muxOutConnector[19] = fifoOut[33][2];
              muxOutConnector[20] = fifoOut[34][2];
              muxOutConnector[21] = fifoOut[35][2];
              muxOutConnector[22] = fifoOut[36][2];
              muxOutConnector[23] = fifoOut[37][2];
              muxOutConnector[24] = fifoOut[38][2];
              muxOutConnector[25] = fifoOut[39][2];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[35][11];
              muxOutConnector[28] = fifoOut[36][11];
              muxOutConnector[29] = fifoOut[37][11];
              muxOutConnector[30] = fifoOut[38][11];
              muxOutConnector[31] = fifoOut[39][11];
              muxOutConnector[32] = fifoOut[40][11];
              muxOutConnector[33] = fifoOut[41][11];
              muxOutConnector[34] = fifoOut[42][11];
              muxOutConnector[35] = fifoOut[43][11];
              muxOutConnector[36] = fifoOut[44][11];
              muxOutConnector[37] = fifoOut[45][11];
              muxOutConnector[38] = fifoOut[46][11];
              muxOutConnector[39] = fifoOut[47][11];
              muxOutConnector[40] = fifoOut[48][11];
              muxOutConnector[41] = fifoOut[49][11];
              muxOutConnector[42] = fifoOut[50][11];
              muxOutConnector[43] = fifoOut[51][11];
              muxOutConnector[44] = fifoOut[26][10];
              muxOutConnector[45] = fifoOut[27][10];
              muxOutConnector[46] = fifoOut[28][10];
              muxOutConnector[47] = fifoOut[29][10];
              muxOutConnector[48] = fifoOut[30][10];
              muxOutConnector[49] = fifoOut[31][10];
              muxOutConnector[50] = fifoOut[32][10];
              muxOutConnector[51] = fifoOut[33][10];
       end
       7: begin
              muxOutConnector[0] = fifoOut[40][3];
              muxOutConnector[1] = fifoOut[41][3];
              muxOutConnector[2] = fifoOut[42][3];
              muxOutConnector[3] = fifoOut[43][3];
              muxOutConnector[4] = fifoOut[44][3];
              muxOutConnector[5] = fifoOut[45][3];
              muxOutConnector[6] = fifoOut[46][3];
              muxOutConnector[7] = fifoOut[47][3];
              muxOutConnector[8] = fifoOut[48][3];
              muxOutConnector[9] = fifoOut[49][3];
              muxOutConnector[10] = fifoOut[50][3];
              muxOutConnector[11] = fifoOut[51][3];
              muxOutConnector[12] = fifoOut[26][2];
              muxOutConnector[13] = fifoOut[27][2];
              muxOutConnector[14] = fifoOut[28][2];
              muxOutConnector[15] = fifoOut[29][2];
              muxOutConnector[16] = fifoOut[30][2];
              muxOutConnector[17] = fifoOut[31][2];
              muxOutConnector[18] = fifoOut[32][2];
              muxOutConnector[19] = fifoOut[33][2];
              muxOutConnector[20] = fifoOut[34][2];
              muxOutConnector[21] = fifoOut[35][2];
              muxOutConnector[22] = fifoOut[36][2];
              muxOutConnector[23] = fifoOut[37][2];
              muxOutConnector[24] = fifoOut[38][2];
              muxOutConnector[25] = fifoOut[39][2];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[35][11];
              muxOutConnector[28] = fifoOut[36][11];
              muxOutConnector[29] = fifoOut[37][11];
              muxOutConnector[30] = fifoOut[38][11];
              muxOutConnector[31] = fifoOut[39][11];
              muxOutConnector[32] = fifoOut[40][11];
              muxOutConnector[33] = fifoOut[41][11];
              muxOutConnector[34] = fifoOut[42][11];
              muxOutConnector[35] = fifoOut[43][11];
              muxOutConnector[36] = fifoOut[44][11];
              muxOutConnector[37] = fifoOut[45][11];
              muxOutConnector[38] = fifoOut[46][11];
              muxOutConnector[39] = fifoOut[47][11];
              muxOutConnector[40] = fifoOut[48][11];
              muxOutConnector[41] = fifoOut[49][11];
              muxOutConnector[42] = fifoOut[50][11];
              muxOutConnector[43] = fifoOut[51][11];
              muxOutConnector[44] = fifoOut[26][10];
              muxOutConnector[45] = fifoOut[27][10];
              muxOutConnector[46] = fifoOut[28][10];
              muxOutConnector[47] = fifoOut[29][10];
              muxOutConnector[48] = fifoOut[30][10];
              muxOutConnector[49] = fifoOut[31][10];
              muxOutConnector[50] = fifoOut[32][10];
              muxOutConnector[51] = fifoOut[33][10];
       end
       8: begin
              muxOutConnector[0] = fifoOut[40][3];
              muxOutConnector[1] = fifoOut[41][3];
              muxOutConnector[2] = fifoOut[42][3];
              muxOutConnector[3] = fifoOut[43][3];
              muxOutConnector[4] = fifoOut[44][3];
              muxOutConnector[5] = fifoOut[45][3];
              muxOutConnector[6] = fifoOut[46][3];
              muxOutConnector[7] = fifoOut[47][3];
              muxOutConnector[8] = fifoOut[48][3];
              muxOutConnector[9] = fifoOut[49][3];
              muxOutConnector[10] = fifoOut[50][3];
              muxOutConnector[11] = fifoOut[51][3];
              muxOutConnector[12] = fifoOut[26][2];
              muxOutConnector[13] = fifoOut[27][2];
              muxOutConnector[14] = fifoOut[28][2];
              muxOutConnector[15] = fifoOut[29][2];
              muxOutConnector[16] = fifoOut[30][2];
              muxOutConnector[17] = fifoOut[31][2];
              muxOutConnector[18] = fifoOut[32][2];
              muxOutConnector[19] = fifoOut[33][2];
              muxOutConnector[20] = fifoOut[34][2];
              muxOutConnector[21] = fifoOut[0][7];
              muxOutConnector[22] = fifoOut[1][7];
              muxOutConnector[23] = fifoOut[2][7];
              muxOutConnector[24] = fifoOut[3][7];
              muxOutConnector[25] = fifoOut[4][7];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[35][11];
              muxOutConnector[28] = fifoOut[36][11];
              muxOutConnector[29] = fifoOut[37][11];
              muxOutConnector[30] = fifoOut[38][11];
              muxOutConnector[31] = fifoOut[39][11];
              muxOutConnector[32] = fifoOut[40][11];
              muxOutConnector[33] = fifoOut[41][11];
              muxOutConnector[34] = fifoOut[42][11];
              muxOutConnector[35] = fifoOut[43][11];
              muxOutConnector[36] = fifoOut[44][11];
              muxOutConnector[37] = fifoOut[45][11];
              muxOutConnector[38] = fifoOut[46][11];
              muxOutConnector[39] = fifoOut[47][11];
              muxOutConnector[40] = fifoOut[48][11];
              muxOutConnector[41] = fifoOut[49][11];
              muxOutConnector[42] = fifoOut[50][11];
              muxOutConnector[43] = fifoOut[51][11];
              muxOutConnector[44] = fifoOut[26][10];
              muxOutConnector[45] = fifoOut[27][10];
              muxOutConnector[46] = fifoOut[28][10];
              muxOutConnector[47] = fifoOut[29][10];
              muxOutConnector[48] = fifoOut[30][10];
              muxOutConnector[49] = fifoOut[31][10];
              muxOutConnector[50] = fifoOut[32][10];
              muxOutConnector[51] = fifoOut[33][10];
       end
       9: begin
              muxOutConnector[0] = fifoOut[5][8];
              muxOutConnector[1] = fifoOut[6][8];
              muxOutConnector[2] = fifoOut[7][8];
              muxOutConnector[3] = fifoOut[8][8];
              muxOutConnector[4] = fifoOut[9][8];
              muxOutConnector[5] = fifoOut[10][8];
              muxOutConnector[6] = fifoOut[11][8];
              muxOutConnector[7] = fifoOut[12][8];
              muxOutConnector[8] = fifoOut[13][8];
              muxOutConnector[9] = fifoOut[14][8];
              muxOutConnector[10] = fifoOut[15][8];
              muxOutConnector[11] = fifoOut[16][8];
              muxOutConnector[12] = fifoOut[17][8];
              muxOutConnector[13] = fifoOut[18][8];
              muxOutConnector[14] = fifoOut[19][8];
              muxOutConnector[15] = fifoOut[20][8];
              muxOutConnector[16] = fifoOut[21][8];
              muxOutConnector[17] = fifoOut[22][8];
              muxOutConnector[18] = fifoOut[23][8];
              muxOutConnector[19] = fifoOut[24][8];
              muxOutConnector[20] = fifoOut[25][8];
              muxOutConnector[21] = fifoOut[0][7];
              muxOutConnector[22] = fifoOut[1][7];
              muxOutConnector[23] = fifoOut[2][7];
              muxOutConnector[24] = fifoOut[3][7];
              muxOutConnector[25] = fifoOut[4][7];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[35][11];
              muxOutConnector[28] = fifoOut[36][11];
              muxOutConnector[29] = fifoOut[37][11];
              muxOutConnector[30] = fifoOut[38][11];
              muxOutConnector[31] = fifoOut[39][11];
              muxOutConnector[32] = fifoOut[40][11];
              muxOutConnector[33] = fifoOut[41][11];
              muxOutConnector[34] = fifoOut[42][11];
              muxOutConnector[35] = fifoOut[43][11];
              muxOutConnector[36] = fifoOut[44][11];
              muxOutConnector[37] = fifoOut[45][11];
              muxOutConnector[38] = fifoOut[46][11];
              muxOutConnector[39] = fifoOut[47][11];
              muxOutConnector[40] = fifoOut[48][11];
              muxOutConnector[41] = fifoOut[49][11];
              muxOutConnector[42] = fifoOut[50][11];
              muxOutConnector[43] = fifoOut[51][11];
              muxOutConnector[44] = fifoOut[26][10];
              muxOutConnector[45] = fifoOut[27][10];
              muxOutConnector[46] = fifoOut[28][10];
              muxOutConnector[47] = fifoOut[29][10];
              muxOutConnector[48] = fifoOut[30][10];
              muxOutConnector[49] = fifoOut[31][10];
              muxOutConnector[50] = fifoOut[32][10];
              muxOutConnector[51] = fifoOut[33][10];
       end
       10: begin
              muxOutConnector[0] = fifoOut[5][8];
              muxOutConnector[1] = fifoOut[6][8];
              muxOutConnector[2] = fifoOut[7][8];
              muxOutConnector[3] = fifoOut[8][8];
              muxOutConnector[4] = fifoOut[9][8];
              muxOutConnector[5] = fifoOut[10][8];
              muxOutConnector[6] = fifoOut[11][8];
              muxOutConnector[7] = fifoOut[12][8];
              muxOutConnector[8] = fifoOut[13][8];
              muxOutConnector[9] = fifoOut[14][8];
              muxOutConnector[10] = fifoOut[15][8];
              muxOutConnector[11] = fifoOut[16][8];
              muxOutConnector[12] = fifoOut[17][8];
              muxOutConnector[13] = fifoOut[18][8];
              muxOutConnector[14] = fifoOut[19][8];
              muxOutConnector[15] = fifoOut[20][8];
              muxOutConnector[16] = fifoOut[21][8];
              muxOutConnector[17] = fifoOut[22][8];
              muxOutConnector[18] = fifoOut[23][8];
              muxOutConnector[19] = fifoOut[24][8];
              muxOutConnector[20] = fifoOut[25][8];
              muxOutConnector[21] = fifoOut[0][7];
              muxOutConnector[22] = fifoOut[1][7];
              muxOutConnector[23] = fifoOut[2][7];
              muxOutConnector[24] = fifoOut[3][7];
              muxOutConnector[25] = fifoOut[4][7];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[35][11];
              muxOutConnector[28] = fifoOut[36][11];
              muxOutConnector[29] = fifoOut[37][11];
              muxOutConnector[30] = fifoOut[38][11];
              muxOutConnector[31] = fifoOut[39][11];
              muxOutConnector[32] = fifoOut[40][11];
              muxOutConnector[33] = fifoOut[41][11];
              muxOutConnector[34] = fifoOut[42][11];
              muxOutConnector[35] = fifoOut[43][11];
              muxOutConnector[36] = fifoOut[44][11];
              muxOutConnector[37] = fifoOut[45][11];
              muxOutConnector[38] = fifoOut[46][11];
              muxOutConnector[39] = fifoOut[47][11];
              muxOutConnector[40] = fifoOut[48][11];
              muxOutConnector[41] = fifoOut[49][11];
              muxOutConnector[42] = fifoOut[50][11];
              muxOutConnector[43] = fifoOut[51][11];
              muxOutConnector[44] = fifoOut[26][10];
              muxOutConnector[45] = fifoOut[27][10];
              muxOutConnector[46] = fifoOut[28][10];
              muxOutConnector[47] = fifoOut[29][10];
              muxOutConnector[48] = fifoOut[30][10];
              muxOutConnector[49] = fifoOut[31][10];
              muxOutConnector[50] = fifoOut[32][10];
              muxOutConnector[51] = fifoOut[33][10];
       end
       11: begin
              muxOutConnector[0] = fifoOut[5][8];
              muxOutConnector[1] = fifoOut[6][8];
              muxOutConnector[2] = fifoOut[7][8];
              muxOutConnector[3] = fifoOut[8][8];
              muxOutConnector[4] = fifoOut[9][8];
              muxOutConnector[5] = fifoOut[10][8];
              muxOutConnector[6] = fifoOut[11][8];
              muxOutConnector[7] = fifoOut[12][8];
              muxOutConnector[8] = fifoOut[13][8];
              muxOutConnector[9] = fifoOut[14][8];
              muxOutConnector[10] = fifoOut[15][8];
              muxOutConnector[11] = fifoOut[16][8];
              muxOutConnector[12] = fifoOut[17][8];
              muxOutConnector[13] = fifoOut[18][8];
              muxOutConnector[14] = fifoOut[19][8];
              muxOutConnector[15] = fifoOut[20][8];
              muxOutConnector[16] = fifoOut[21][8];
              muxOutConnector[17] = fifoOut[22][8];
              muxOutConnector[18] = fifoOut[23][8];
              muxOutConnector[19] = fifoOut[24][8];
              muxOutConnector[20] = fifoOut[25][8];
              muxOutConnector[21] = fifoOut[0][7];
              muxOutConnector[22] = fifoOut[1][7];
              muxOutConnector[23] = fifoOut[2][7];
              muxOutConnector[24] = fifoOut[3][7];
              muxOutConnector[25] = fifoOut[4][7];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[35][11];
              muxOutConnector[28] = fifoOut[36][11];
              muxOutConnector[29] = fifoOut[37][11];
              muxOutConnector[30] = fifoOut[38][11];
              muxOutConnector[31] = fifoOut[39][11];
              muxOutConnector[32] = fifoOut[40][11];
              muxOutConnector[33] = fifoOut[41][11];
              muxOutConnector[34] = fifoOut[42][11];
              muxOutConnector[35] = fifoOut[8][1];
              muxOutConnector[36] = fifoOut[9][1];
              muxOutConnector[37] = fifoOut[10][1];
              muxOutConnector[38] = fifoOut[11][1];
              muxOutConnector[39] = fifoOut[12][1];
              muxOutConnector[40] = fifoOut[13][1];
              muxOutConnector[41] = fifoOut[14][1];
              muxOutConnector[42] = fifoOut[15][1];
              muxOutConnector[43] = fifoOut[16][1];
              muxOutConnector[44] = fifoOut[17][1];
              muxOutConnector[45] = fifoOut[18][1];
              muxOutConnector[46] = fifoOut[19][1];
              muxOutConnector[47] = fifoOut[20][1];
              muxOutConnector[48] = fifoOut[21][1];
              muxOutConnector[49] = fifoOut[22][1];
              muxOutConnector[50] = fifoOut[23][1];
              muxOutConnector[51] = fifoOut[24][1];
       end
       12: begin
              muxOutConnector[0] = fifoOut[5][8];
              muxOutConnector[1] = fifoOut[6][8];
              muxOutConnector[2] = fifoOut[7][8];
              muxOutConnector[3] = fifoOut[8][8];
              muxOutConnector[4] = fifoOut[9][8];
              muxOutConnector[5] = fifoOut[10][8];
              muxOutConnector[6] = fifoOut[11][8];
              muxOutConnector[7] = fifoOut[12][8];
              muxOutConnector[8] = fifoOut[13][8];
              muxOutConnector[9] = fifoOut[14][8];
              muxOutConnector[10] = fifoOut[15][8];
              muxOutConnector[11] = fifoOut[16][8];
              muxOutConnector[12] = fifoOut[17][8];
              muxOutConnector[13] = fifoOut[18][8];
              muxOutConnector[14] = fifoOut[19][8];
              muxOutConnector[15] = fifoOut[20][8];
              muxOutConnector[16] = fifoOut[21][8];
              muxOutConnector[17] = fifoOut[22][8];
              muxOutConnector[18] = fifoOut[23][8];
              muxOutConnector[19] = fifoOut[24][8];
              muxOutConnector[20] = fifoOut[25][8];
              muxOutConnector[21] = fifoOut[0][7];
              muxOutConnector[22] = fifoOut[1][7];
              muxOutConnector[23] = fifoOut[2][7];
              muxOutConnector[24] = fifoOut[3][7];
              muxOutConnector[25] = fifoOut[4][7];
              muxOutConnector[26] = fifoOut[25][2];
              muxOutConnector[27] = fifoOut[0][1];
              muxOutConnector[28] = fifoOut[1][1];
              muxOutConnector[29] = fifoOut[2][1];
              muxOutConnector[30] = fifoOut[3][1];
              muxOutConnector[31] = fifoOut[4][1];
              muxOutConnector[32] = fifoOut[5][1];
              muxOutConnector[33] = fifoOut[6][1];
              muxOutConnector[34] = fifoOut[7][1];
              muxOutConnector[35] = fifoOut[8][1];
              muxOutConnector[36] = fifoOut[9][1];
              muxOutConnector[37] = fifoOut[10][1];
              muxOutConnector[38] = fifoOut[11][1];
              muxOutConnector[39] = fifoOut[12][1];
              muxOutConnector[40] = fifoOut[13][1];
              muxOutConnector[41] = fifoOut[14][1];
              muxOutConnector[42] = fifoOut[15][1];
              muxOutConnector[43] = fifoOut[16][1];
              muxOutConnector[44] = fifoOut[17][1];
              muxOutConnector[45] = fifoOut[18][1];
              muxOutConnector[46] = fifoOut[19][1];
              muxOutConnector[47] = fifoOut[20][1];
              muxOutConnector[48] = fifoOut[21][1];
              muxOutConnector[49] = fifoOut[22][1];
              muxOutConnector[50] = fifoOut[23][1];
              muxOutConnector[51] = fifoOut[24][1];
       end
       13: begin
              muxOutConnector[0] = fifoOut[5][8];
              muxOutConnector[1] = fifoOut[6][8];
              muxOutConnector[2] = fifoOut[7][8];
              muxOutConnector[3] = fifoOut[8][8];
              muxOutConnector[4] = fifoOut[9][8];
              muxOutConnector[5] = fifoOut[10][8];
              muxOutConnector[6] = fifoOut[11][8];
              muxOutConnector[7] = fifoOut[12][8];
              muxOutConnector[8] = fifoOut[13][8];
              muxOutConnector[9] = fifoOut[14][8];
              muxOutConnector[10] = fifoOut[15][8];
              muxOutConnector[11] = fifoOut[16][8];
              muxOutConnector[12] = fifoOut[17][8];
              muxOutConnector[13] = fifoOut[18][8];
              muxOutConnector[14] = fifoOut[19][8];
              muxOutConnector[15] = fifoOut[20][8];
              muxOutConnector[16] = fifoOut[21][8];
              muxOutConnector[17] = fifoOut[22][8];
              muxOutConnector[18] = fifoOut[23][8];
              muxOutConnector[19] = fifoOut[24][8];
              muxOutConnector[20] = fifoOut[25][8];
              muxOutConnector[21] = fifoOut[0][7];
              muxOutConnector[22] = fifoOut[1][7];
              muxOutConnector[23] = fifoOut[2][7];
              muxOutConnector[24] = fifoOut[3][7];
              muxOutConnector[25] = fifoOut[4][7];
              muxOutConnector[26] = fifoOut[25][2];
              muxOutConnector[27] = fifoOut[0][1];
              muxOutConnector[28] = fifoOut[1][1];
              muxOutConnector[29] = fifoOut[2][1];
              muxOutConnector[30] = fifoOut[3][1];
              muxOutConnector[31] = fifoOut[4][1];
              muxOutConnector[32] = fifoOut[5][1];
              muxOutConnector[33] = fifoOut[6][1];
              muxOutConnector[34] = fifoOut[7][1];
              muxOutConnector[35] = fifoOut[8][1];
              muxOutConnector[36] = fifoOut[9][1];
              muxOutConnector[37] = fifoOut[10][1];
              muxOutConnector[38] = fifoOut[11][1];
              muxOutConnector[39] = fifoOut[12][1];
              muxOutConnector[40] = fifoOut[13][1];
              muxOutConnector[41] = fifoOut[14][1];
              muxOutConnector[42] = fifoOut[15][1];
              muxOutConnector[43] = fifoOut[16][1];
              muxOutConnector[44] = fifoOut[17][1];
              muxOutConnector[45] = fifoOut[18][1];
              muxOutConnector[46] = fifoOut[19][1];
              muxOutConnector[47] = fifoOut[20][1];
              muxOutConnector[48] = fifoOut[21][1];
              muxOutConnector[49] = fifoOut[22][1];
              muxOutConnector[50] = fifoOut[23][1];
              muxOutConnector[51] = fifoOut[24][1];
       end
       14: begin
              muxOutConnector[0] = fifoOut[5][8];
              muxOutConnector[1] = fifoOut[6][8];
              muxOutConnector[2] = fifoOut[7][8];
              muxOutConnector[3] = fifoOut[8][8];
              muxOutConnector[4] = fifoOut[9][8];
              muxOutConnector[5] = fifoOut[10][8];
              muxOutConnector[6] = fifoOut[11][8];
              muxOutConnector[7] = fifoOut[12][8];
              muxOutConnector[8] = fifoOut[13][8];
              muxOutConnector[9] = fifoOut[14][8];
              muxOutConnector[10] = fifoOut[15][8];
              muxOutConnector[11] = fifoOut[16][8];
              muxOutConnector[12] = fifoOut[17][8];
              muxOutConnector[13] = fifoOut[18][8];
              muxOutConnector[14] = fifoOut[19][8];
              muxOutConnector[15] = fifoOut[20][8];
              muxOutConnector[16] = fifoOut[21][8];
              muxOutConnector[17] = fifoOut[22][8];
              muxOutConnector[18] = fifoOut[23][8];
              muxOutConnector[19] = fifoOut[24][8];
              muxOutConnector[20] = fifoOut[25][8];
              muxOutConnector[21] = fifoOut[0][7];
              muxOutConnector[22] = fifoOut[1][7];
              muxOutConnector[23] = fifoOut[2][7];
              muxOutConnector[24] = fifoOut[3][7];
              muxOutConnector[25] = fifoOut[4][7];
              muxOutConnector[26] = fifoOut[25][2];
              muxOutConnector[27] = fifoOut[0][1];
              muxOutConnector[28] = fifoOut[1][1];
              muxOutConnector[29] = fifoOut[2][1];
              muxOutConnector[30] = fifoOut[3][1];
              muxOutConnector[31] = fifoOut[4][1];
              muxOutConnector[32] = fifoOut[5][1];
              muxOutConnector[33] = fifoOut[6][1];
              muxOutConnector[34] = fifoOut[7][1];
              muxOutConnector[35] = fifoOut[8][1];
              muxOutConnector[36] = fifoOut[9][1];
              muxOutConnector[37] = fifoOut[10][1];
              muxOutConnector[38] = fifoOut[11][1];
              muxOutConnector[39] = fifoOut[12][1];
              muxOutConnector[40] = fifoOut[13][1];
              muxOutConnector[41] = fifoOut[14][1];
              muxOutConnector[42] = fifoOut[15][1];
              muxOutConnector[43] = fifoOut[16][1];
              muxOutConnector[44] = fifoOut[17][1];
              muxOutConnector[45] = fifoOut[18][1];
              muxOutConnector[46] = fifoOut[19][1];
              muxOutConnector[47] = fifoOut[20][1];
              muxOutConnector[48] = fifoOut[21][1];
              muxOutConnector[49] = fifoOut[22][1];
              muxOutConnector[50] = fifoOut[23][1];
              muxOutConnector[51] = fifoOut[24][1];
       end
       15: begin
              muxOutConnector[0] = fifoOut[5][8];
              muxOutConnector[1] = fifoOut[6][8];
              muxOutConnector[2] = fifoOut[7][8];
              muxOutConnector[3] = fifoOut[8][8];
              muxOutConnector[4] = fifoOut[9][8];
              muxOutConnector[5] = fifoOut[10][8];
              muxOutConnector[6] = fifoOut[11][8];
              muxOutConnector[7] = fifoOut[12][8];
              muxOutConnector[8] = fifoOut[13][8];
              muxOutConnector[9] = fifoOut[14][8];
              muxOutConnector[10] = fifoOut[15][8];
              muxOutConnector[11] = fifoOut[16][8];
              muxOutConnector[12] = fifoOut[17][8];
              muxOutConnector[13] = fifoOut[18][8];
              muxOutConnector[14] = fifoOut[19][8];
              muxOutConnector[15] = fifoOut[20][8];
              muxOutConnector[16] = fifoOut[21][8];
              muxOutConnector[17] = fifoOut[22][8];
              muxOutConnector[18] = fifoOut[23][8];
              muxOutConnector[19] = fifoOut[24][8];
              muxOutConnector[20] = fifoOut[25][8];
              muxOutConnector[21] = fifoOut[0][7];
              muxOutConnector[22] = fifoOut[1][7];
              muxOutConnector[23] = fifoOut[2][7];
              muxOutConnector[24] = fifoOut[3][7];
              muxOutConnector[25] = fifoOut[4][7];
              muxOutConnector[26] = fifoOut[25][2];
              muxOutConnector[27] = fifoOut[0][1];
              muxOutConnector[28] = fifoOut[1][1];
              muxOutConnector[29] = fifoOut[2][1];
              muxOutConnector[30] = fifoOut[3][1];
              muxOutConnector[31] = fifoOut[4][1];
              muxOutConnector[32] = fifoOut[5][1];
              muxOutConnector[33] = fifoOut[6][1];
              muxOutConnector[34] = fifoOut[7][1];
              muxOutConnector[35] = fifoOut[8][1];
              muxOutConnector[36] = fifoOut[9][1];
              muxOutConnector[37] = fifoOut[10][1];
              muxOutConnector[38] = fifoOut[11][1];
              muxOutConnector[39] = fifoOut[12][1];
              muxOutConnector[40] = fifoOut[13][1];
              muxOutConnector[41] = fifoOut[14][1];
              muxOutConnector[42] = fifoOut[15][1];
              muxOutConnector[43] = fifoOut[16][1];
              muxOutConnector[44] = fifoOut[17][1];
              muxOutConnector[45] = fifoOut[18][1];
              muxOutConnector[46] = fifoOut[19][1];
              muxOutConnector[47] = fifoOut[20][1];
              muxOutConnector[48] = fifoOut[21][1];
              muxOutConnector[49] = fifoOut[22][1];
              muxOutConnector[50] = fifoOut[23][1];
              muxOutConnector[51] = fifoOut[24][1];
       end
       16: begin
              muxOutConnector[0] = fifoOut[5][8];
              muxOutConnector[1] = fifoOut[6][8];
              muxOutConnector[2] = fifoOut[7][8];
              muxOutConnector[3] = fifoOut[8][8];
              muxOutConnector[4] = fifoOut[9][8];
              muxOutConnector[5] = fifoOut[10][8];
              muxOutConnector[6] = fifoOut[11][8];
              muxOutConnector[7] = fifoOut[12][8];
              muxOutConnector[8] = fifoOut[13][8];
              muxOutConnector[9] = fifoOut[14][8];
              muxOutConnector[10] = fifoOut[15][8];
              muxOutConnector[11] = fifoOut[16][8];
              muxOutConnector[12] = fifoOut[17][8];
              muxOutConnector[13] = fifoOut[18][8];
              muxOutConnector[14] = fifoOut[19][8];
              muxOutConnector[15] = fifoOut[20][8];
              muxOutConnector[16] = fifoOut[21][8];
              muxOutConnector[17] = fifoOut[22][8];
              muxOutConnector[18] = fifoOut[23][8];
              muxOutConnector[19] = fifoOut[24][8];
              muxOutConnector[20] = fifoOut[25][8];
              muxOutConnector[21] = fifoOut[0][7];
              muxOutConnector[22] = fifoOut[1][7];
              muxOutConnector[23] = fifoOut[2][7];
              muxOutConnector[24] = fifoOut[3][7];
              muxOutConnector[25] = fifoOut[4][7];
              muxOutConnector[26] = fifoOut[25][2];
              muxOutConnector[27] = fifoOut[0][1];
              muxOutConnector[28] = fifoOut[1][1];
              muxOutConnector[29] = fifoOut[2][1];
              muxOutConnector[30] = fifoOut[3][1];
              muxOutConnector[31] = fifoOut[4][1];
              muxOutConnector[32] = fifoOut[5][1];
              muxOutConnector[33] = fifoOut[6][1];
              muxOutConnector[34] = fifoOut[7][1];
              muxOutConnector[35] = fifoOut[8][1];
              muxOutConnector[36] = fifoOut[9][1];
              muxOutConnector[37] = fifoOut[10][1];
              muxOutConnector[38] = fifoOut[11][1];
              muxOutConnector[39] = fifoOut[12][1];
              muxOutConnector[40] = fifoOut[13][1];
              muxOutConnector[41] = fifoOut[14][1];
              muxOutConnector[42] = fifoOut[15][1];
              muxOutConnector[43] = fifoOut[16][1];
              muxOutConnector[44] = fifoOut[35][0];
              muxOutConnector[45] = fifoOut[36][0];
              muxOutConnector[46] = fifoOut[37][0];
              muxOutConnector[47] = fifoOut[38][0];
              muxOutConnector[48] = fifoOut[39][0];
              muxOutConnector[49] = fifoOut[40][0];
              muxOutConnector[50] = fifoOut[41][0];
              muxOutConnector[51] = fifoOut[42][0];
       end
       17: begin
              muxOutConnector[0] = fifoOut[5][8];
              muxOutConnector[1] = fifoOut[6][8];
              muxOutConnector[2] = fifoOut[7][8];
              muxOutConnector[3] = fifoOut[8][8];
              muxOutConnector[4] = fifoOut[9][8];
              muxOutConnector[5] = fifoOut[10][8];
              muxOutConnector[6] = fifoOut[11][8];
              muxOutConnector[7] = fifoOut[12][8];
              muxOutConnector[8] = fifoOut[13][8];
              muxOutConnector[9] = fifoOut[14][8];
              muxOutConnector[10] = fifoOut[15][8];
              muxOutConnector[11] = fifoOut[16][8];
              muxOutConnector[12] = fifoOut[17][8];
              muxOutConnector[13] = fifoOut[18][8];
              muxOutConnector[14] = fifoOut[19][8];
              muxOutConnector[15] = fifoOut[20][8];
              muxOutConnector[16] = fifoOut[21][8];
              muxOutConnector[17] = fifoOut[22][8];
              muxOutConnector[18] = fifoOut[23][8];
              muxOutConnector[19] = fifoOut[24][8];
              muxOutConnector[20] = fifoOut[25][8];
              muxOutConnector[21] = fifoOut[0][7];
              muxOutConnector[22] = fifoOut[1][7];
              muxOutConnector[23] = fifoOut[2][7];
              muxOutConnector[24] = fifoOut[3][7];
              muxOutConnector[25] = fifoOut[4][7];
              muxOutConnector[26] = fifoOut[43][1];
              muxOutConnector[27] = fifoOut[44][1];
              muxOutConnector[28] = fifoOut[45][1];
              muxOutConnector[29] = fifoOut[46][1];
              muxOutConnector[30] = fifoOut[47][1];
              muxOutConnector[31] = fifoOut[48][1];
              muxOutConnector[32] = fifoOut[49][1];
              muxOutConnector[33] = fifoOut[50][1];
              muxOutConnector[34] = fifoOut[51][1];
              muxOutConnector[35] = fifoOut[26][0];
              muxOutConnector[36] = fifoOut[27][0];
              muxOutConnector[37] = fifoOut[28][0];
              muxOutConnector[38] = fifoOut[29][0];
              muxOutConnector[39] = fifoOut[30][0];
              muxOutConnector[40] = fifoOut[31][0];
              muxOutConnector[41] = fifoOut[32][0];
              muxOutConnector[42] = fifoOut[33][0];
              muxOutConnector[43] = fifoOut[34][0];
              muxOutConnector[44] = fifoOut[35][0];
              muxOutConnector[45] = fifoOut[36][0];
              muxOutConnector[46] = fifoOut[37][0];
              muxOutConnector[47] = fifoOut[38][0];
              muxOutConnector[48] = fifoOut[39][0];
              muxOutConnector[49] = fifoOut[40][0];
              muxOutConnector[50] = fifoOut[41][0];
              muxOutConnector[51] = fifoOut[42][0];
       end
       18: begin
              muxOutConnector[0] = fifoOut[5][8];
              muxOutConnector[1] = fifoOut[6][8];
              muxOutConnector[2] = fifoOut[7][8];
              muxOutConnector[3] = fifoOut[8][8];
              muxOutConnector[4] = fifoOut[9][8];
              muxOutConnector[5] = fifoOut[10][8];
              muxOutConnector[6] = fifoOut[11][8];
              muxOutConnector[7] = fifoOut[12][8];
              muxOutConnector[8] = fifoOut[13][8];
              muxOutConnector[9] = fifoOut[14][8];
              muxOutConnector[10] = fifoOut[15][8];
              muxOutConnector[11] = fifoOut[16][8];
              muxOutConnector[12] = fifoOut[17][8];
              muxOutConnector[13] = fifoOut[18][8];
              muxOutConnector[14] = fifoOut[19][8];
              muxOutConnector[15] = fifoOut[20][8];
              muxOutConnector[16] = fifoOut[21][8];
              muxOutConnector[17] = fifoOut[22][8];
              muxOutConnector[18] = fifoOut[23][8];
              muxOutConnector[19] = fifoOut[24][8];
              muxOutConnector[20] = fifoOut[25][8];
              muxOutConnector[21] = fifoOut[0][7];
              muxOutConnector[22] = fifoOut[1][7];
              muxOutConnector[23] = fifoOut[2][7];
              muxOutConnector[24] = fifoOut[3][7];
              muxOutConnector[25] = fifoOut[4][7];
              muxOutConnector[26] = fifoOut[43][1];
              muxOutConnector[27] = fifoOut[44][1];
              muxOutConnector[28] = fifoOut[45][1];
              muxOutConnector[29] = fifoOut[46][1];
              muxOutConnector[30] = fifoOut[47][1];
              muxOutConnector[31] = fifoOut[48][1];
              muxOutConnector[32] = fifoOut[49][1];
              muxOutConnector[33] = fifoOut[50][1];
              muxOutConnector[34] = fifoOut[51][1];
              muxOutConnector[35] = fifoOut[26][0];
              muxOutConnector[36] = fifoOut[27][0];
              muxOutConnector[37] = fifoOut[28][0];
              muxOutConnector[38] = fifoOut[29][0];
              muxOutConnector[39] = fifoOut[30][0];
              muxOutConnector[40] = fifoOut[31][0];
              muxOutConnector[41] = fifoOut[32][0];
              muxOutConnector[42] = fifoOut[33][0];
              muxOutConnector[43] = fifoOut[34][0];
              muxOutConnector[44] = fifoOut[35][0];
              muxOutConnector[45] = fifoOut[36][0];
              muxOutConnector[46] = fifoOut[37][0];
              muxOutConnector[47] = fifoOut[38][0];
              muxOutConnector[48] = fifoOut[39][0];
              muxOutConnector[49] = fifoOut[40][0];
              muxOutConnector[50] = fifoOut[41][0];
              muxOutConnector[51] = fifoOut[42][0];
       end
       19: begin
              muxOutConnector[0] = fifoOut[5][8];
              muxOutConnector[1] = fifoOut[6][8];
              muxOutConnector[2] = fifoOut[7][8];
              muxOutConnector[3] = fifoOut[8][8];
              muxOutConnector[4] = fifoOut[9][8];
              muxOutConnector[5] = fifoOut[10][8];
              muxOutConnector[6] = fifoOut[11][8];
              muxOutConnector[7] = fifoOut[12][8];
              muxOutConnector[8] = fifoOut[13][8];
              muxOutConnector[9] = fifoOut[14][8];
              muxOutConnector[10] = fifoOut[15][8];
              muxOutConnector[11] = fifoOut[16][8];
              muxOutConnector[12] = fifoOut[17][8];
              muxOutConnector[13] = fifoOut[18][8];
              muxOutConnector[14] = fifoOut[19][8];
              muxOutConnector[15] = fifoOut[20][8];
              muxOutConnector[16] = fifoOut[21][8];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[43][1];
              muxOutConnector[27] = fifoOut[44][1];
              muxOutConnector[28] = fifoOut[45][1];
              muxOutConnector[29] = fifoOut[46][1];
              muxOutConnector[30] = fifoOut[47][1];
              muxOutConnector[31] = fifoOut[48][1];
              muxOutConnector[32] = fifoOut[49][1];
              muxOutConnector[33] = fifoOut[50][1];
              muxOutConnector[34] = fifoOut[51][1];
              muxOutConnector[35] = fifoOut[26][0];
              muxOutConnector[36] = fifoOut[27][0];
              muxOutConnector[37] = fifoOut[28][0];
              muxOutConnector[38] = fifoOut[29][0];
              muxOutConnector[39] = fifoOut[30][0];
              muxOutConnector[40] = fifoOut[31][0];
              muxOutConnector[41] = fifoOut[32][0];
              muxOutConnector[42] = fifoOut[33][0];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
