`timescale 1ns / 1ps
module LMem1To0_511_circ6_yesshift_nounload_scripted(
        muxOut,
        ly0In,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 14;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            fifoOut[i][0] <= ly0InConnector[i];
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[21][2];
              muxOutConnector[1] = fifoOut[22][2];
              muxOutConnector[2] = fifoOut[23][2];
              muxOutConnector[3] = fifoOut[24][2];
              muxOutConnector[4] = fifoOut[25][2];
              muxOutConnector[5] = fifoOut[0][1];
              muxOutConnector[6] = fifoOut[1][1];
              muxOutConnector[7] = fifoOut[2][1];
              muxOutConnector[8] = fifoOut[3][1];
              muxOutConnector[9] = fifoOut[4][1];
              muxOutConnector[10] = fifoOut[5][1];
              muxOutConnector[11] = fifoOut[6][1];
              muxOutConnector[12] = fifoOut[7][1];
              muxOutConnector[13] = fifoOut[8][1];
              muxOutConnector[14] = fifoOut[9][1];
              muxOutConnector[15] = fifoOut[10][1];
              muxOutConnector[16] = fifoOut[11][1];
              muxOutConnector[17] = fifoOut[12][1];
              muxOutConnector[18] = fifoOut[13][1];
              muxOutConnector[19] = fifoOut[14][1];
              muxOutConnector[20] = fifoOut[15][1];
              muxOutConnector[21] = fifoOut[16][1];
              muxOutConnector[22] = fifoOut[17][1];
              muxOutConnector[23] = fifoOut[18][1];
              muxOutConnector[24] = fifoOut[19][1];
              muxOutConnector[25] = fifoOut[20][1];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
       end
       1: begin
              muxOutConnector[0] = fifoOut[21][2];
              muxOutConnector[1] = fifoOut[22][2];
              muxOutConnector[2] = fifoOut[23][2];
              muxOutConnector[3] = fifoOut[24][2];
              muxOutConnector[4] = fifoOut[25][2];
              muxOutConnector[5] = fifoOut[0][1];
              muxOutConnector[6] = fifoOut[1][1];
              muxOutConnector[7] = fifoOut[2][1];
              muxOutConnector[8] = fifoOut[3][1];
              muxOutConnector[9] = fifoOut[4][1];
              muxOutConnector[10] = fifoOut[5][1];
              muxOutConnector[11] = fifoOut[6][1];
              muxOutConnector[12] = fifoOut[7][1];
              muxOutConnector[13] = fifoOut[8][1];
              muxOutConnector[14] = fifoOut[9][1];
              muxOutConnector[15] = fifoOut[10][1];
              muxOutConnector[16] = fifoOut[11][1];
              muxOutConnector[17] = fifoOut[12][1];
              muxOutConnector[18] = fifoOut[13][1];
              muxOutConnector[19] = fifoOut[14][1];
              muxOutConnector[20] = fifoOut[15][1];
              muxOutConnector[21] = fifoOut[16][1];
              muxOutConnector[22] = fifoOut[33][0];
              muxOutConnector[23] = fifoOut[34][0];
              muxOutConnector[24] = fifoOut[35][0];
              muxOutConnector[25] = fifoOut[36][0];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
       end
       2: begin
              muxOutConnector[0] = fifoOut[37][1];
              muxOutConnector[1] = fifoOut[38][1];
              muxOutConnector[2] = fifoOut[39][1];
              muxOutConnector[3] = fifoOut[40][1];
              muxOutConnector[4] = fifoOut[41][1];
              muxOutConnector[5] = fifoOut[42][1];
              muxOutConnector[6] = fifoOut[43][1];
              muxOutConnector[7] = fifoOut[44][1];
              muxOutConnector[8] = fifoOut[45][1];
              muxOutConnector[9] = fifoOut[46][1];
              muxOutConnector[10] = fifoOut[47][1];
              muxOutConnector[11] = fifoOut[48][1];
              muxOutConnector[12] = fifoOut[49][1];
              muxOutConnector[13] = fifoOut[50][1];
              muxOutConnector[14] = fifoOut[51][1];
              muxOutConnector[15] = fifoOut[26][0];
              muxOutConnector[16] = fifoOut[27][0];
              muxOutConnector[17] = fifoOut[28][0];
              muxOutConnector[18] = fifoOut[29][0];
              muxOutConnector[19] = fifoOut[30][0];
              muxOutConnector[20] = fifoOut[31][0];
              muxOutConnector[21] = fifoOut[32][0];
              muxOutConnector[22] = fifoOut[33][0];
              muxOutConnector[23] = fifoOut[34][0];
              muxOutConnector[24] = fifoOut[35][0];
              muxOutConnector[25] = fifoOut[36][0];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
       end
       3: begin
              muxOutConnector[0] = fifoOut[37][1];
              muxOutConnector[1] = fifoOut[38][1];
              muxOutConnector[2] = fifoOut[39][1];
              muxOutConnector[3] = fifoOut[40][1];
              muxOutConnector[4] = fifoOut[41][1];
              muxOutConnector[5] = fifoOut[42][1];
              muxOutConnector[6] = fifoOut[43][1];
              muxOutConnector[7] = fifoOut[44][1];
              muxOutConnector[8] = fifoOut[45][1];
              muxOutConnector[9] = fifoOut[46][1];
              muxOutConnector[10] = fifoOut[47][1];
              muxOutConnector[11] = fifoOut[48][1];
              muxOutConnector[12] = fifoOut[49][1];
              muxOutConnector[13] = fifoOut[50][1];
              muxOutConnector[14] = fifoOut[51][1];
              muxOutConnector[15] = fifoOut[26][0];
              muxOutConnector[16] = fifoOut[27][0];
              muxOutConnector[17] = fifoOut[28][0];
              muxOutConnector[18] = fifoOut[29][0];
              muxOutConnector[19] = fifoOut[30][0];
              muxOutConnector[20] = fifoOut[31][0];
              muxOutConnector[21] = fifoOut[32][0];
              muxOutConnector[22] = fifoOut[33][0];
              muxOutConnector[23] = fifoOut[34][0];
              muxOutConnector[24] = fifoOut[35][0];
              muxOutConnector[25] = fifoOut[36][0];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
       end
       4: begin
              muxOutConnector[0] = fifoOut[37][1];
              muxOutConnector[1] = fifoOut[38][1];
              muxOutConnector[2] = fifoOut[39][1];
              muxOutConnector[3] = fifoOut[40][1];
              muxOutConnector[4] = fifoOut[41][1];
              muxOutConnector[5] = fifoOut[42][1];
              muxOutConnector[6] = fifoOut[43][1];
              muxOutConnector[7] = fifoOut[44][1];
              muxOutConnector[8] = fifoOut[45][1];
              muxOutConnector[9] = fifoOut[46][1];
              muxOutConnector[10] = fifoOut[47][1];
              muxOutConnector[11] = fifoOut[48][1];
              muxOutConnector[12] = fifoOut[49][1];
              muxOutConnector[13] = fifoOut[50][1];
              muxOutConnector[14] = fifoOut[51][1];
              muxOutConnector[15] = fifoOut[26][0];
              muxOutConnector[16] = fifoOut[27][0];
              muxOutConnector[17] = fifoOut[28][0];
              muxOutConnector[18] = fifoOut[29][0];
              muxOutConnector[19] = fifoOut[30][0];
              muxOutConnector[20] = fifoOut[31][0];
              muxOutConnector[21] = fifoOut[32][0];
              muxOutConnector[22] = fifoOut[33][0];
              muxOutConnector[23] = fifoOut[34][0];
              muxOutConnector[24] = fifoOut[35][0];
              muxOutConnector[25] = fifoOut[36][0];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
       end
       5: begin
              muxOutConnector[0] = fifoOut[37][1];
              muxOutConnector[1] = fifoOut[38][1];
              muxOutConnector[2] = fifoOut[39][1];
              muxOutConnector[3] = fifoOut[40][1];
              muxOutConnector[4] = fifoOut[41][1];
              muxOutConnector[5] = fifoOut[42][1];
              muxOutConnector[6] = fifoOut[43][1];
              muxOutConnector[7] = fifoOut[44][1];
              muxOutConnector[8] = fifoOut[45][1];
              muxOutConnector[9] = fifoOut[46][1];
              muxOutConnector[10] = fifoOut[47][1];
              muxOutConnector[11] = fifoOut[48][1];
              muxOutConnector[12] = fifoOut[49][1];
              muxOutConnector[13] = fifoOut[50][1];
              muxOutConnector[14] = fifoOut[51][1];
              muxOutConnector[15] = fifoOut[26][0];
              muxOutConnector[16] = fifoOut[27][0];
              muxOutConnector[17] = fifoOut[28][0];
              muxOutConnector[18] = fifoOut[29][0];
              muxOutConnector[19] = fifoOut[30][0];
              muxOutConnector[20] = fifoOut[31][0];
              muxOutConnector[21] = fifoOut[32][0];
              muxOutConnector[22] = fifoOut[33][0];
              muxOutConnector[23] = fifoOut[34][0];
              muxOutConnector[24] = fifoOut[35][0];
              muxOutConnector[25] = fifoOut[36][0];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
       end
       6: begin
              muxOutConnector[0] = fifoOut[37][1];
              muxOutConnector[1] = fifoOut[38][1];
              muxOutConnector[2] = fifoOut[39][1];
              muxOutConnector[3] = fifoOut[40][1];
              muxOutConnector[4] = fifoOut[41][1];
              muxOutConnector[5] = fifoOut[42][1];
              muxOutConnector[6] = fifoOut[43][1];
              muxOutConnector[7] = fifoOut[44][1];
              muxOutConnector[8] = fifoOut[45][1];
              muxOutConnector[9] = fifoOut[46][1];
              muxOutConnector[10] = fifoOut[47][1];
              muxOutConnector[11] = fifoOut[48][1];
              muxOutConnector[12] = fifoOut[49][1];
              muxOutConnector[13] = fifoOut[50][1];
              muxOutConnector[14] = fifoOut[51][1];
              muxOutConnector[15] = fifoOut[26][0];
              muxOutConnector[16] = fifoOut[27][0];
              muxOutConnector[17] = fifoOut[28][0];
              muxOutConnector[18] = fifoOut[29][0];
              muxOutConnector[19] = fifoOut[30][0];
              muxOutConnector[20] = fifoOut[31][0];
              muxOutConnector[21] = fifoOut[32][0];
              muxOutConnector[22] = fifoOut[33][0];
              muxOutConnector[23] = fifoOut[34][0];
              muxOutConnector[24] = fifoOut[35][0];
              muxOutConnector[25] = fifoOut[36][0];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
       end
       7: begin
              muxOutConnector[0] = fifoOut[37][1];
              muxOutConnector[1] = fifoOut[38][1];
              muxOutConnector[2] = fifoOut[39][1];
              muxOutConnector[3] = fifoOut[40][1];
              muxOutConnector[4] = fifoOut[41][1];
              muxOutConnector[5] = fifoOut[42][1];
              muxOutConnector[6] = fifoOut[43][1];
              muxOutConnector[7] = fifoOut[44][1];
              muxOutConnector[8] = fifoOut[45][1];
              muxOutConnector[9] = fifoOut[46][1];
              muxOutConnector[10] = fifoOut[47][1];
              muxOutConnector[11] = fifoOut[48][1];
              muxOutConnector[12] = fifoOut[49][1];
              muxOutConnector[13] = fifoOut[50][1];
              muxOutConnector[14] = fifoOut[51][1];
              muxOutConnector[15] = fifoOut[26][0];
              muxOutConnector[16] = fifoOut[27][0];
              muxOutConnector[17] = fifoOut[28][0];
              muxOutConnector[18] = fifoOut[29][0];
              muxOutConnector[19] = fifoOut[30][0];
              muxOutConnector[20] = fifoOut[31][0];
              muxOutConnector[21] = fifoOut[32][0];
              muxOutConnector[22] = fifoOut[0][6];
              muxOutConnector[23] = fifoOut[1][6];
              muxOutConnector[24] = fifoOut[2][6];
              muxOutConnector[25] = fifoOut[3][6];
              muxOutConnector[26] = fifoOut[17][8];
              muxOutConnector[27] = fifoOut[18][8];
              muxOutConnector[28] = fifoOut[19][8];
              muxOutConnector[29] = fifoOut[20][8];
              muxOutConnector[30] = fifoOut[21][8];
              muxOutConnector[31] = fifoOut[22][8];
              muxOutConnector[32] = fifoOut[23][8];
              muxOutConnector[33] = fifoOut[24][8];
              muxOutConnector[34] = fifoOut[25][8];
              muxOutConnector[35] = fifoOut[0][7];
              muxOutConnector[36] = fifoOut[1][7];
              muxOutConnector[37] = fifoOut[2][7];
              muxOutConnector[38] = fifoOut[3][7];
              muxOutConnector[39] = fifoOut[4][7];
              muxOutConnector[40] = fifoOut[5][7];
              muxOutConnector[41] = fifoOut[6][7];
              muxOutConnector[42] = fifoOut[7][7];
              muxOutConnector[43] = fifoOut[8][7];
              muxOutConnector[44] = fifoOut[9][7];
              muxOutConnector[45] = fifoOut[10][7];
              muxOutConnector[46] = fifoOut[11][7];
              muxOutConnector[47] = fifoOut[12][7];
              muxOutConnector[48] = fifoOut[13][7];
              muxOutConnector[49] = fifoOut[14][7];
              muxOutConnector[50] = fifoOut[15][7];
              muxOutConnector[51] = fifoOut[16][7];
       end
       8: begin
              muxOutConnector[0] = fifoOut[4][7];
              muxOutConnector[1] = fifoOut[5][7];
              muxOutConnector[2] = fifoOut[6][7];
              muxOutConnector[3] = fifoOut[7][7];
              muxOutConnector[4] = fifoOut[8][7];
              muxOutConnector[5] = fifoOut[9][7];
              muxOutConnector[6] = fifoOut[10][7];
              muxOutConnector[7] = fifoOut[11][7];
              muxOutConnector[8] = fifoOut[12][7];
              muxOutConnector[9] = fifoOut[13][7];
              muxOutConnector[10] = fifoOut[14][7];
              muxOutConnector[11] = fifoOut[15][7];
              muxOutConnector[12] = fifoOut[16][7];
              muxOutConnector[13] = fifoOut[17][7];
              muxOutConnector[14] = fifoOut[18][7];
              muxOutConnector[15] = fifoOut[19][7];
              muxOutConnector[16] = fifoOut[20][7];
              muxOutConnector[17] = fifoOut[21][7];
              muxOutConnector[18] = fifoOut[22][7];
              muxOutConnector[19] = fifoOut[23][7];
              muxOutConnector[20] = fifoOut[24][7];
              muxOutConnector[21] = fifoOut[25][7];
              muxOutConnector[22] = fifoOut[0][6];
              muxOutConnector[23] = fifoOut[1][6];
              muxOutConnector[24] = fifoOut[2][6];
              muxOutConnector[25] = fifoOut[3][6];
              muxOutConnector[26] = fifoOut[33][7];
              muxOutConnector[27] = fifoOut[34][7];
              muxOutConnector[28] = fifoOut[35][7];
              muxOutConnector[29] = fifoOut[36][7];
              muxOutConnector[30] = fifoOut[37][7];
              muxOutConnector[31] = fifoOut[38][7];
              muxOutConnector[32] = fifoOut[39][7];
              muxOutConnector[33] = fifoOut[40][7];
              muxOutConnector[34] = fifoOut[41][7];
              muxOutConnector[35] = fifoOut[42][7];
              muxOutConnector[36] = fifoOut[43][7];
              muxOutConnector[37] = fifoOut[44][7];
              muxOutConnector[38] = fifoOut[45][7];
              muxOutConnector[39] = fifoOut[46][7];
              muxOutConnector[40] = fifoOut[47][7];
              muxOutConnector[41] = fifoOut[48][7];
              muxOutConnector[42] = fifoOut[49][7];
              muxOutConnector[43] = fifoOut[50][7];
              muxOutConnector[44] = fifoOut[51][7];
              muxOutConnector[45] = fifoOut[26][6];
              muxOutConnector[46] = fifoOut[27][6];
              muxOutConnector[47] = fifoOut[28][6];
              muxOutConnector[48] = fifoOut[29][6];
              muxOutConnector[49] = fifoOut[30][6];
              muxOutConnector[50] = fifoOut[31][6];
              muxOutConnector[51] = fifoOut[32][6];
       end
       9: begin
              muxOutConnector[0] = fifoOut[4][7];
              muxOutConnector[1] = fifoOut[5][7];
              muxOutConnector[2] = fifoOut[6][7];
              muxOutConnector[3] = fifoOut[7][7];
              muxOutConnector[4] = fifoOut[8][7];
              muxOutConnector[5] = fifoOut[9][7];
              muxOutConnector[6] = fifoOut[10][7];
              muxOutConnector[7] = fifoOut[11][7];
              muxOutConnector[8] = fifoOut[12][7];
              muxOutConnector[9] = fifoOut[13][7];
              muxOutConnector[10] = fifoOut[14][7];
              muxOutConnector[11] = fifoOut[15][7];
              muxOutConnector[12] = fifoOut[16][7];
              muxOutConnector[13] = fifoOut[17][7];
              muxOutConnector[14] = fifoOut[18][7];
              muxOutConnector[15] = fifoOut[19][7];
              muxOutConnector[16] = fifoOut[20][7];
              muxOutConnector[17] = fifoOut[21][7];
              muxOutConnector[18] = fifoOut[22][7];
              muxOutConnector[19] = fifoOut[23][7];
              muxOutConnector[20] = fifoOut[24][7];
              muxOutConnector[21] = fifoOut[25][7];
              muxOutConnector[22] = fifoOut[0][6];
              muxOutConnector[23] = fifoOut[1][6];
              muxOutConnector[24] = fifoOut[2][6];
              muxOutConnector[25] = fifoOut[3][6];
              muxOutConnector[26] = fifoOut[33][7];
              muxOutConnector[27] = fifoOut[34][7];
              muxOutConnector[28] = fifoOut[35][7];
              muxOutConnector[29] = fifoOut[36][7];
              muxOutConnector[30] = fifoOut[37][7];
              muxOutConnector[31] = fifoOut[38][7];
              muxOutConnector[32] = fifoOut[39][7];
              muxOutConnector[33] = fifoOut[40][7];
              muxOutConnector[34] = fifoOut[41][7];
              muxOutConnector[35] = fifoOut[42][7];
              muxOutConnector[36] = fifoOut[43][7];
              muxOutConnector[37] = fifoOut[44][7];
              muxOutConnector[38] = fifoOut[45][7];
              muxOutConnector[39] = fifoOut[46][7];
              muxOutConnector[40] = fifoOut[47][7];
              muxOutConnector[41] = fifoOut[48][7];
              muxOutConnector[42] = fifoOut[49][7];
              muxOutConnector[43] = fifoOut[50][7];
              muxOutConnector[44] = fifoOut[51][7];
              muxOutConnector[45] = fifoOut[26][6];
              muxOutConnector[46] = fifoOut[27][6];
              muxOutConnector[47] = fifoOut[28][6];
              muxOutConnector[48] = fifoOut[29][6];
              muxOutConnector[49] = fifoOut[30][6];
              muxOutConnector[50] = fifoOut[31][6];
              muxOutConnector[51] = fifoOut[32][6];
       end
       10: begin
              muxOutConnector[0] = fifoOut[4][7];
              muxOutConnector[1] = fifoOut[5][7];
              muxOutConnector[2] = fifoOut[6][7];
              muxOutConnector[3] = fifoOut[7][7];
              muxOutConnector[4] = fifoOut[8][7];
              muxOutConnector[5] = fifoOut[9][7];
              muxOutConnector[6] = fifoOut[10][7];
              muxOutConnector[7] = fifoOut[11][7];
              muxOutConnector[8] = fifoOut[12][7];
              muxOutConnector[9] = fifoOut[13][7];
              muxOutConnector[10] = fifoOut[14][7];
              muxOutConnector[11] = fifoOut[15][7];
              muxOutConnector[12] = fifoOut[16][7];
              muxOutConnector[13] = fifoOut[17][7];
              muxOutConnector[14] = fifoOut[18][7];
              muxOutConnector[15] = fifoOut[19][7];
              muxOutConnector[16] = fifoOut[20][7];
              muxOutConnector[17] = fifoOut[21][7];
              muxOutConnector[18] = fifoOut[22][7];
              muxOutConnector[19] = fifoOut[23][7];
              muxOutConnector[20] = fifoOut[24][7];
              muxOutConnector[21] = fifoOut[25][7];
              muxOutConnector[22] = fifoOut[0][6];
              muxOutConnector[23] = fifoOut[1][6];
              muxOutConnector[24] = fifoOut[2][6];
              muxOutConnector[25] = fifoOut[3][6];
              muxOutConnector[26] = fifoOut[33][7];
              muxOutConnector[27] = fifoOut[34][7];
              muxOutConnector[28] = fifoOut[35][7];
              muxOutConnector[29] = fifoOut[36][7];
              muxOutConnector[30] = fifoOut[37][7];
              muxOutConnector[31] = fifoOut[38][7];
              muxOutConnector[32] = fifoOut[39][7];
              muxOutConnector[33] = fifoOut[40][7];
              muxOutConnector[34] = fifoOut[41][7];
              muxOutConnector[35] = fifoOut[42][7];
              muxOutConnector[36] = fifoOut[43][7];
              muxOutConnector[37] = fifoOut[44][7];
              muxOutConnector[38] = fifoOut[45][7];
              muxOutConnector[39] = fifoOut[46][7];
              muxOutConnector[40] = fifoOut[47][7];
              muxOutConnector[41] = fifoOut[48][7];
              muxOutConnector[42] = fifoOut[49][7];
              muxOutConnector[43] = fifoOut[50][7];
              muxOutConnector[44] = fifoOut[51][7];
              muxOutConnector[45] = fifoOut[26][6];
              muxOutConnector[46] = fifoOut[27][6];
              muxOutConnector[47] = fifoOut[28][6];
              muxOutConnector[48] = fifoOut[29][6];
              muxOutConnector[49] = fifoOut[30][6];
              muxOutConnector[50] = fifoOut[31][6];
              muxOutConnector[51] = fifoOut[32][6];
       end
       11: begin
              muxOutConnector[0] = fifoOut[4][7];
              muxOutConnector[1] = fifoOut[5][7];
              muxOutConnector[2] = fifoOut[6][7];
              muxOutConnector[3] = fifoOut[7][7];
              muxOutConnector[4] = fifoOut[8][7];
              muxOutConnector[5] = fifoOut[9][7];
              muxOutConnector[6] = fifoOut[10][7];
              muxOutConnector[7] = fifoOut[11][7];
              muxOutConnector[8] = fifoOut[12][7];
              muxOutConnector[9] = fifoOut[13][7];
              muxOutConnector[10] = fifoOut[14][7];
              muxOutConnector[11] = fifoOut[15][7];
              muxOutConnector[12] = fifoOut[16][7];
              muxOutConnector[13] = fifoOut[17][7];
              muxOutConnector[14] = fifoOut[18][7];
              muxOutConnector[15] = fifoOut[19][7];
              muxOutConnector[16] = fifoOut[20][7];
              muxOutConnector[17] = fifoOut[21][7];
              muxOutConnector[18] = fifoOut[22][7];
              muxOutConnector[19] = fifoOut[23][7];
              muxOutConnector[20] = fifoOut[24][7];
              muxOutConnector[21] = fifoOut[25][7];
              muxOutConnector[22] = fifoOut[0][6];
              muxOutConnector[23] = fifoOut[1][6];
              muxOutConnector[24] = fifoOut[2][6];
              muxOutConnector[25] = fifoOut[3][6];
              muxOutConnector[26] = fifoOut[33][7];
              muxOutConnector[27] = fifoOut[34][7];
              muxOutConnector[28] = fifoOut[35][7];
              muxOutConnector[29] = fifoOut[36][7];
              muxOutConnector[30] = fifoOut[37][7];
              muxOutConnector[31] = fifoOut[38][7];
              muxOutConnector[32] = fifoOut[39][7];
              muxOutConnector[33] = fifoOut[40][7];
              muxOutConnector[34] = fifoOut[41][7];
              muxOutConnector[35] = fifoOut[42][7];
              muxOutConnector[36] = fifoOut[43][7];
              muxOutConnector[37] = fifoOut[44][7];
              muxOutConnector[38] = fifoOut[45][7];
              muxOutConnector[39] = fifoOut[46][7];
              muxOutConnector[40] = fifoOut[47][7];
              muxOutConnector[41] = fifoOut[48][7];
              muxOutConnector[42] = fifoOut[49][7];
              muxOutConnector[43] = fifoOut[50][7];
              muxOutConnector[44] = fifoOut[51][7];
              muxOutConnector[45] = fifoOut[26][6];
              muxOutConnector[46] = fifoOut[27][6];
              muxOutConnector[47] = fifoOut[28][6];
              muxOutConnector[48] = fifoOut[29][6];
              muxOutConnector[49] = fifoOut[30][6];
              muxOutConnector[50] = fifoOut[31][6];
              muxOutConnector[51] = fifoOut[32][6];
       end
       12: begin
              muxOutConnector[0] = fifoOut[4][7];
              muxOutConnector[1] = fifoOut[5][7];
              muxOutConnector[2] = fifoOut[6][7];
              muxOutConnector[3] = fifoOut[7][7];
              muxOutConnector[4] = fifoOut[8][7];
              muxOutConnector[5] = fifoOut[9][7];
              muxOutConnector[6] = fifoOut[10][7];
              muxOutConnector[7] = fifoOut[11][7];
              muxOutConnector[8] = fifoOut[12][7];
              muxOutConnector[9] = fifoOut[13][7];
              muxOutConnector[10] = fifoOut[14][7];
              muxOutConnector[11] = fifoOut[15][7];
              muxOutConnector[12] = fifoOut[16][7];
              muxOutConnector[13] = fifoOut[17][7];
              muxOutConnector[14] = fifoOut[18][7];
              muxOutConnector[15] = fifoOut[19][7];
              muxOutConnector[16] = fifoOut[20][7];
              muxOutConnector[17] = fifoOut[21][7];
              muxOutConnector[18] = fifoOut[22][7];
              muxOutConnector[19] = fifoOut[23][7];
              muxOutConnector[20] = fifoOut[24][7];
              muxOutConnector[21] = fifoOut[25][7];
              muxOutConnector[22] = fifoOut[0][6];
              muxOutConnector[23] = fifoOut[1][6];
              muxOutConnector[24] = fifoOut[2][6];
              muxOutConnector[25] = fifoOut[3][6];
              muxOutConnector[26] = fifoOut[33][7];
              muxOutConnector[27] = fifoOut[34][7];
              muxOutConnector[28] = fifoOut[35][7];
              muxOutConnector[29] = fifoOut[36][7];
              muxOutConnector[30] = fifoOut[37][7];
              muxOutConnector[31] = fifoOut[38][7];
              muxOutConnector[32] = fifoOut[39][7];
              muxOutConnector[33] = fifoOut[40][7];
              muxOutConnector[34] = fifoOut[41][7];
              muxOutConnector[35] = fifoOut[42][7];
              muxOutConnector[36] = fifoOut[43][7];
              muxOutConnector[37] = fifoOut[44][7];
              muxOutConnector[38] = fifoOut[45][7];
              muxOutConnector[39] = fifoOut[46][7];
              muxOutConnector[40] = fifoOut[47][7];
              muxOutConnector[41] = fifoOut[48][7];
              muxOutConnector[42] = fifoOut[49][7];
              muxOutConnector[43] = fifoOut[50][7];
              muxOutConnector[44] = fifoOut[51][7];
              muxOutConnector[45] = fifoOut[26][6];
              muxOutConnector[46] = fifoOut[27][6];
              muxOutConnector[47] = fifoOut[28][6];
              muxOutConnector[48] = fifoOut[29][6];
              muxOutConnector[49] = fifoOut[30][6];
              muxOutConnector[50] = fifoOut[31][6];
              muxOutConnector[51] = fifoOut[32][6];
       end
       13: begin
              muxOutConnector[0] = fifoOut[4][7];
              muxOutConnector[1] = fifoOut[5][7];
              muxOutConnector[2] = fifoOut[6][7];
              muxOutConnector[3] = fifoOut[7][7];
              muxOutConnector[4] = fifoOut[8][7];
              muxOutConnector[5] = fifoOut[9][7];
              muxOutConnector[6] = fifoOut[10][7];
              muxOutConnector[7] = fifoOut[11][7];
              muxOutConnector[8] = fifoOut[12][7];
              muxOutConnector[9] = fifoOut[13][7];
              muxOutConnector[10] = fifoOut[14][7];
              muxOutConnector[11] = fifoOut[15][7];
              muxOutConnector[12] = fifoOut[16][7];
              muxOutConnector[13] = fifoOut[17][7];
              muxOutConnector[14] = fifoOut[18][7];
              muxOutConnector[15] = fifoOut[19][7];
              muxOutConnector[16] = fifoOut[20][7];
              muxOutConnector[17] = fifoOut[21][7];
              muxOutConnector[18] = fifoOut[22][7];
              muxOutConnector[19] = fifoOut[23][7];
              muxOutConnector[20] = fifoOut[24][7];
              muxOutConnector[21] = fifoOut[25][7];
              muxOutConnector[22] = fifoOut[0][6];
              muxOutConnector[23] = fifoOut[1][6];
              muxOutConnector[24] = fifoOut[2][6];
              muxOutConnector[25] = fifoOut[3][6];
              muxOutConnector[26] = fifoOut[33][7];
              muxOutConnector[27] = fifoOut[34][7];
              muxOutConnector[28] = fifoOut[35][7];
              muxOutConnector[29] = fifoOut[36][7];
              muxOutConnector[30] = fifoOut[37][7];
              muxOutConnector[31] = fifoOut[38][7];
              muxOutConnector[32] = fifoOut[39][7];
              muxOutConnector[33] = fifoOut[40][7];
              muxOutConnector[34] = fifoOut[41][7];
              muxOutConnector[35] = fifoOut[42][7];
              muxOutConnector[36] = fifoOut[43][7];
              muxOutConnector[37] = fifoOut[44][7];
              muxOutConnector[38] = fifoOut[45][7];
              muxOutConnector[39] = fifoOut[46][7];
              muxOutConnector[40] = fifoOut[47][7];
              muxOutConnector[41] = fifoOut[48][7];
              muxOutConnector[42] = fifoOut[49][7];
              muxOutConnector[43] = fifoOut[50][7];
              muxOutConnector[44] = fifoOut[51][7];
              muxOutConnector[45] = fifoOut[26][6];
              muxOutConnector[46] = fifoOut[27][6];
              muxOutConnector[47] = fifoOut[28][6];
              muxOutConnector[48] = fifoOut[29][6];
              muxOutConnector[49] = fifoOut[30][6];
              muxOutConnector[50] = fifoOut[31][6];
              muxOutConnector[51] = fifoOut[32][6];
       end
       14: begin
              muxOutConnector[0] = fifoOut[4][7];
              muxOutConnector[1] = fifoOut[5][7];
              muxOutConnector[2] = fifoOut[6][7];
              muxOutConnector[3] = fifoOut[7][7];
              muxOutConnector[4] = fifoOut[8][7];
              muxOutConnector[5] = fifoOut[9][7];
              muxOutConnector[6] = fifoOut[10][7];
              muxOutConnector[7] = fifoOut[11][7];
              muxOutConnector[8] = fifoOut[12][7];
              muxOutConnector[9] = fifoOut[13][7];
              muxOutConnector[10] = fifoOut[14][7];
              muxOutConnector[11] = fifoOut[15][7];
              muxOutConnector[12] = fifoOut[16][7];
              muxOutConnector[13] = fifoOut[17][7];
              muxOutConnector[14] = fifoOut[18][7];
              muxOutConnector[15] = fifoOut[19][7];
              muxOutConnector[16] = fifoOut[20][7];
              muxOutConnector[17] = fifoOut[21][7];
              muxOutConnector[18] = fifoOut[22][7];
              muxOutConnector[19] = fifoOut[23][7];
              muxOutConnector[20] = fifoOut[24][7];
              muxOutConnector[21] = fifoOut[25][7];
              muxOutConnector[22] = fifoOut[0][6];
              muxOutConnector[23] = fifoOut[1][6];
              muxOutConnector[24] = fifoOut[2][6];
              muxOutConnector[25] = fifoOut[3][6];
              muxOutConnector[26] = fifoOut[0][13];
              muxOutConnector[27] = fifoOut[1][13];
              muxOutConnector[28] = fifoOut[2][13];
              muxOutConnector[29] = fifoOut[3][13];
              muxOutConnector[30] = fifoOut[4][13];
              muxOutConnector[31] = fifoOut[5][13];
              muxOutConnector[32] = fifoOut[6][13];
              muxOutConnector[33] = fifoOut[7][13];
              muxOutConnector[34] = fifoOut[8][13];
              muxOutConnector[35] = fifoOut[9][13];
              muxOutConnector[36] = fifoOut[10][13];
              muxOutConnector[37] = fifoOut[11][13];
              muxOutConnector[38] = fifoOut[12][13];
              muxOutConnector[39] = fifoOut[13][13];
              muxOutConnector[40] = fifoOut[14][13];
              muxOutConnector[41] = fifoOut[15][13];
              muxOutConnector[42] = fifoOut[16][13];
              muxOutConnector[43] = fifoOut[17][13];
              muxOutConnector[44] = fifoOut[18][13];
              muxOutConnector[45] = fifoOut[19][13];
              muxOutConnector[46] = fifoOut[20][13];
              muxOutConnector[47] = fifoOut[21][13];
              muxOutConnector[48] = fifoOut[22][13];
              muxOutConnector[49] = fifoOut[23][13];
              muxOutConnector[50] = fifoOut[24][13];
              muxOutConnector[51] = fifoOut[25][13];
       end
       15: begin
              muxOutConnector[0] = fifoOut[4][7];
              muxOutConnector[1] = fifoOut[5][7];
              muxOutConnector[2] = fifoOut[6][7];
              muxOutConnector[3] = fifoOut[7][7];
              muxOutConnector[4] = fifoOut[8][7];
              muxOutConnector[5] = fifoOut[9][7];
              muxOutConnector[6] = fifoOut[10][7];
              muxOutConnector[7] = fifoOut[11][7];
              muxOutConnector[8] = fifoOut[12][7];
              muxOutConnector[9] = fifoOut[13][7];
              muxOutConnector[10] = fifoOut[14][7];
              muxOutConnector[11] = fifoOut[15][7];
              muxOutConnector[12] = fifoOut[16][7];
              muxOutConnector[13] = fifoOut[17][7];
              muxOutConnector[14] = fifoOut[18][7];
              muxOutConnector[15] = fifoOut[19][7];
              muxOutConnector[16] = fifoOut[20][7];
              muxOutConnector[17] = fifoOut[21][7];
              muxOutConnector[18] = fifoOut[22][7];
              muxOutConnector[19] = fifoOut[23][7];
              muxOutConnector[20] = fifoOut[24][7];
              muxOutConnector[21] = fifoOut[25][7];
              muxOutConnector[22] = fifoOut[0][6];
              muxOutConnector[23] = fifoOut[1][6];
              muxOutConnector[24] = fifoOut[2][6];
              muxOutConnector[25] = fifoOut[3][6];
              muxOutConnector[26] = fifoOut[0][13];
              muxOutConnector[27] = fifoOut[1][13];
              muxOutConnector[28] = fifoOut[2][13];
              muxOutConnector[29] = fifoOut[3][13];
              muxOutConnector[30] = fifoOut[4][13];
              muxOutConnector[31] = fifoOut[5][13];
              muxOutConnector[32] = fifoOut[6][13];
              muxOutConnector[33] = fifoOut[7][13];
              muxOutConnector[34] = fifoOut[8][13];
              muxOutConnector[35] = fifoOut[9][13];
              muxOutConnector[36] = fifoOut[10][13];
              muxOutConnector[37] = fifoOut[11][13];
              muxOutConnector[38] = fifoOut[12][13];
              muxOutConnector[39] = fifoOut[13][13];
              muxOutConnector[40] = fifoOut[14][13];
              muxOutConnector[41] = fifoOut[15][13];
              muxOutConnector[42] = fifoOut[16][13];
              muxOutConnector[43] = fifoOut[17][13];
              muxOutConnector[44] = fifoOut[18][13];
              muxOutConnector[45] = fifoOut[19][13];
              muxOutConnector[46] = fifoOut[20][13];
              muxOutConnector[47] = fifoOut[21][13];
              muxOutConnector[48] = fifoOut[22][13];
              muxOutConnector[49] = fifoOut[23][13];
              muxOutConnector[50] = fifoOut[24][13];
              muxOutConnector[51] = fifoOut[25][13];
       end
       16: begin
              muxOutConnector[0] = fifoOut[4][7];
              muxOutConnector[1] = fifoOut[5][7];
              muxOutConnector[2] = fifoOut[6][7];
              muxOutConnector[3] = fifoOut[7][7];
              muxOutConnector[4] = fifoOut[8][7];
              muxOutConnector[5] = fifoOut[9][7];
              muxOutConnector[6] = fifoOut[10][7];
              muxOutConnector[7] = fifoOut[11][7];
              muxOutConnector[8] = fifoOut[12][7];
              muxOutConnector[9] = fifoOut[13][7];
              muxOutConnector[10] = fifoOut[14][7];
              muxOutConnector[11] = fifoOut[15][7];
              muxOutConnector[12] = fifoOut[16][7];
              muxOutConnector[13] = fifoOut[17][7];
              muxOutConnector[14] = fifoOut[18][7];
              muxOutConnector[15] = fifoOut[19][7];
              muxOutConnector[16] = fifoOut[20][7];
              muxOutConnector[17] = fifoOut[21][7];
              muxOutConnector[18] = fifoOut[22][7];
              muxOutConnector[19] = fifoOut[23][7];
              muxOutConnector[20] = fifoOut[24][7];
              muxOutConnector[21] = fifoOut[25][7];
              muxOutConnector[22] = fifoOut[0][6];
              muxOutConnector[23] = fifoOut[1][6];
              muxOutConnector[24] = fifoOut[2][6];
              muxOutConnector[25] = fifoOut[3][6];
              muxOutConnector[26] = fifoOut[0][13];
              muxOutConnector[27] = fifoOut[1][13];
              muxOutConnector[28] = fifoOut[2][13];
              muxOutConnector[29] = fifoOut[3][13];
              muxOutConnector[30] = fifoOut[4][13];
              muxOutConnector[31] = fifoOut[5][13];
              muxOutConnector[32] = fifoOut[6][13];
              muxOutConnector[33] = fifoOut[7][13];
              muxOutConnector[34] = fifoOut[8][13];
              muxOutConnector[35] = fifoOut[9][13];
              muxOutConnector[36] = fifoOut[10][13];
              muxOutConnector[37] = fifoOut[11][13];
              muxOutConnector[38] = fifoOut[12][13];
              muxOutConnector[39] = fifoOut[13][13];
              muxOutConnector[40] = fifoOut[14][13];
              muxOutConnector[41] = fifoOut[15][13];
              muxOutConnector[42] = fifoOut[16][13];
              muxOutConnector[43] = fifoOut[17][13];
              muxOutConnector[44] = fifoOut[18][13];
              muxOutConnector[45] = fifoOut[19][13];
              muxOutConnector[46] = fifoOut[20][13];
              muxOutConnector[47] = fifoOut[21][13];
              muxOutConnector[48] = fifoOut[22][13];
              muxOutConnector[49] = fifoOut[23][13];
              muxOutConnector[50] = fifoOut[24][13];
              muxOutConnector[51] = fifoOut[25][13];
       end
       17: begin
              muxOutConnector[0] = fifoOut[4][7];
              muxOutConnector[1] = fifoOut[5][7];
              muxOutConnector[2] = fifoOut[6][7];
              muxOutConnector[3] = fifoOut[7][7];
              muxOutConnector[4] = fifoOut[8][7];
              muxOutConnector[5] = fifoOut[9][7];
              muxOutConnector[6] = fifoOut[10][7];
              muxOutConnector[7] = fifoOut[11][7];
              muxOutConnector[8] = fifoOut[12][7];
              muxOutConnector[9] = fifoOut[13][7];
              muxOutConnector[10] = fifoOut[14][7];
              muxOutConnector[11] = fifoOut[15][7];
              muxOutConnector[12] = fifoOut[16][7];
              muxOutConnector[13] = fifoOut[17][7];
              muxOutConnector[14] = fifoOut[18][7];
              muxOutConnector[15] = fifoOut[19][7];
              muxOutConnector[16] = fifoOut[20][7];
              muxOutConnector[17] = fifoOut[21][7];
              muxOutConnector[18] = fifoOut[22][7];
              muxOutConnector[19] = fifoOut[23][7];
              muxOutConnector[20] = fifoOut[24][7];
              muxOutConnector[21] = fifoOut[25][7];
              muxOutConnector[22] = fifoOut[0][6];
              muxOutConnector[23] = fifoOut[1][6];
              muxOutConnector[24] = fifoOut[2][6];
              muxOutConnector[25] = fifoOut[3][6];
              muxOutConnector[26] = fifoOut[0][13];
              muxOutConnector[27] = fifoOut[1][13];
              muxOutConnector[28] = fifoOut[2][13];
              muxOutConnector[29] = fifoOut[3][13];
              muxOutConnector[30] = fifoOut[4][13];
              muxOutConnector[31] = fifoOut[5][13];
              muxOutConnector[32] = fifoOut[6][13];
              muxOutConnector[33] = fifoOut[7][13];
              muxOutConnector[34] = fifoOut[8][13];
              muxOutConnector[35] = fifoOut[9][13];
              muxOutConnector[36] = fifoOut[10][13];
              muxOutConnector[37] = fifoOut[11][13];
              muxOutConnector[38] = fifoOut[12][13];
              muxOutConnector[39] = fifoOut[13][13];
              muxOutConnector[40] = fifoOut[14][13];
              muxOutConnector[41] = fifoOut[15][13];
              muxOutConnector[42] = fifoOut[16][13];
              muxOutConnector[43] = fifoOut[17][13];
              muxOutConnector[44] = fifoOut[18][13];
              muxOutConnector[45] = fifoOut[19][13];
              muxOutConnector[46] = fifoOut[20][13];
              muxOutConnector[47] = fifoOut[21][13];
              muxOutConnector[48] = fifoOut[22][13];
              muxOutConnector[49] = fifoOut[23][13];
              muxOutConnector[50] = fifoOut[24][13];
              muxOutConnector[51] = fifoOut[25][13];
       end
       18: begin
              muxOutConnector[0] = fifoOut[4][7];
              muxOutConnector[1] = fifoOut[5][7];
              muxOutConnector[2] = fifoOut[6][7];
              muxOutConnector[3] = fifoOut[7][7];
              muxOutConnector[4] = fifoOut[8][7];
              muxOutConnector[5] = fifoOut[9][7];
              muxOutConnector[6] = fifoOut[10][7];
              muxOutConnector[7] = fifoOut[11][7];
              muxOutConnector[8] = fifoOut[12][7];
              muxOutConnector[9] = fifoOut[13][7];
              muxOutConnector[10] = fifoOut[14][7];
              muxOutConnector[11] = fifoOut[15][7];
              muxOutConnector[12] = fifoOut[16][7];
              muxOutConnector[13] = fifoOut[17][7];
              muxOutConnector[14] = fifoOut[18][7];
              muxOutConnector[15] = fifoOut[19][7];
              muxOutConnector[16] = fifoOut[20][7];
              muxOutConnector[17] = fifoOut[21][7];
              muxOutConnector[18] = fifoOut[22][7];
              muxOutConnector[19] = fifoOut[23][7];
              muxOutConnector[20] = fifoOut[24][7];
              muxOutConnector[21] = fifoOut[25][7];
              muxOutConnector[22] = fifoOut[0][6];
              muxOutConnector[23] = fifoOut[1][6];
              muxOutConnector[24] = fifoOut[2][6];
              muxOutConnector[25] = fifoOut[3][6];
              muxOutConnector[26] = fifoOut[0][13];
              muxOutConnector[27] = fifoOut[1][13];
              muxOutConnector[28] = fifoOut[2][13];
              muxOutConnector[29] = fifoOut[3][13];
              muxOutConnector[30] = fifoOut[4][13];
              muxOutConnector[31] = fifoOut[5][13];
              muxOutConnector[32] = fifoOut[6][13];
              muxOutConnector[33] = fifoOut[7][13];
              muxOutConnector[34] = fifoOut[8][13];
              muxOutConnector[35] = fifoOut[9][13];
              muxOutConnector[36] = fifoOut[10][13];
              muxOutConnector[37] = fifoOut[11][13];
              muxOutConnector[38] = fifoOut[12][13];
              muxOutConnector[39] = fifoOut[13][13];
              muxOutConnector[40] = fifoOut[14][13];
              muxOutConnector[41] = fifoOut[15][13];
              muxOutConnector[42] = fifoOut[16][13];
              muxOutConnector[43] = fifoOut[17][13];
              muxOutConnector[44] = fifoOut[18][13];
              muxOutConnector[45] = fifoOut[19][13];
              muxOutConnector[46] = fifoOut[20][13];
              muxOutConnector[47] = fifoOut[21][13];
              muxOutConnector[48] = fifoOut[22][13];
              muxOutConnector[49] = fifoOut[23][13];
              muxOutConnector[50] = fifoOut[24][13];
              muxOutConnector[51] = fifoOut[25][13];
       end
       19: begin
              muxOutConnector[0] = fifoOut[4][7];
              muxOutConnector[1] = fifoOut[5][7];
              muxOutConnector[2] = fifoOut[6][7];
              muxOutConnector[3] = fifoOut[7][7];
              muxOutConnector[4] = fifoOut[8][7];
              muxOutConnector[5] = fifoOut[9][7];
              muxOutConnector[6] = fifoOut[10][7];
              muxOutConnector[7] = fifoOut[11][7];
              muxOutConnector[8] = fifoOut[12][7];
              muxOutConnector[9] = fifoOut[13][7];
              muxOutConnector[10] = fifoOut[14][7];
              muxOutConnector[11] = fifoOut[15][7];
              muxOutConnector[12] = fifoOut[16][7];
              muxOutConnector[13] = fifoOut[17][7];
              muxOutConnector[14] = fifoOut[18][7];
              muxOutConnector[15] = fifoOut[19][7];
              muxOutConnector[16] = fifoOut[20][7];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[0][13];
              muxOutConnector[27] = fifoOut[1][13];
              muxOutConnector[28] = fifoOut[2][13];
              muxOutConnector[29] = fifoOut[3][13];
              muxOutConnector[30] = fifoOut[4][13];
              muxOutConnector[31] = fifoOut[5][13];
              muxOutConnector[32] = fifoOut[6][13];
              muxOutConnector[33] = fifoOut[7][13];
              muxOutConnector[34] = fifoOut[8][13];
              muxOutConnector[35] = fifoOut[9][13];
              muxOutConnector[36] = fifoOut[10][13];
              muxOutConnector[37] = fifoOut[11][13];
              muxOutConnector[38] = fifoOut[12][13];
              muxOutConnector[39] = fifoOut[13][13];
              muxOutConnector[40] = fifoOut[14][13];
              muxOutConnector[41] = fifoOut[15][13];
              muxOutConnector[42] = fifoOut[16][13];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
