`timescale 1ns / 1ps
module LMem1To0_511_circ1_combined_ys_yu_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        rxIn,
        load_input_en,
        iteration_0_indicator,
        feedback_en,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter r_lower = 32;
parameter c = 17;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input load_input_en;
input iteration_0_indicator;
input [ADDRESSWIDTH-1:0]unloadAddress;
input feedback_en;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input [ r_lower * w - 1 : 0 ] rxIn; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
wire [w-1:0]rxInConnector[r_lower-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

generate
    for (k=0;k<r_lower;k=k+1)begin:assign_rx
        assign rxInConnector[k] = rxIn[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            if(feedback_en)begin
                 fifoOut[i][0] <= fifoOut[i][c-1];
            end
            else if(load_input_en)begin
                 if(i < r_lower)begin
                   fifoOut[i][0] = rxInConnector[i];
                 end
                 else begin
                   fifoOut[i][0] = maxVal;
                 end
            end
            else begin
                 fifoOut[i][0] <= ly0InConnector[i];
            end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
       0: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = fifoOut[17][5][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[18][6][w-1];
              unloadMuxOut[1] = fifoOut[19][6][w-1];
              unloadMuxOut[2] = fifoOut[20][6][w-1];
              unloadMuxOut[3] = fifoOut[21][6][w-1];
              unloadMuxOut[4] = fifoOut[22][6][w-1];
              unloadMuxOut[5] = fifoOut[23][6][w-1];
              unloadMuxOut[6] = fifoOut[24][6][w-1];
              unloadMuxOut[7] = fifoOut[25][6][w-1];
              unloadMuxOut[8] = fifoOut[0][5][w-1];
              unloadMuxOut[9] = fifoOut[1][5][w-1];
              unloadMuxOut[10] = fifoOut[2][5][w-1];
              unloadMuxOut[11] = fifoOut[3][5][w-1];
              unloadMuxOut[12] = fifoOut[4][5][w-1];
              unloadMuxOut[13] = fifoOut[5][5][w-1];
              unloadMuxOut[14] = fifoOut[6][5][w-1];
              unloadMuxOut[15] = fifoOut[7][5][w-1];
              unloadMuxOut[16] = fifoOut[8][5][w-1];
              unloadMuxOut[17] = fifoOut[9][5][w-1];
              unloadMuxOut[18] = fifoOut[10][5][w-1];
              unloadMuxOut[19] = fifoOut[11][5][w-1];
              unloadMuxOut[20] = fifoOut[12][5][w-1];
              unloadMuxOut[21] = fifoOut[13][5][w-1];
              unloadMuxOut[22] = fifoOut[14][5][w-1];
              unloadMuxOut[23] = fifoOut[15][5][w-1];
              unloadMuxOut[24] = fifoOut[16][5][w-1];
              unloadMuxOut[25] = fifoOut[17][5][w-1];
              unloadMuxOut[26] = fifoOut[18][5][w-1];
              unloadMuxOut[27] = fifoOut[19][5][w-1];
              unloadMuxOut[28] = fifoOut[20][5][w-1];
              unloadMuxOut[29] = fifoOut[21][5][w-1];
              unloadMuxOut[30] = fifoOut[22][5][w-1];
              unloadMuxOut[31] = fifoOut[23][5][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[24][6][w-1];
              unloadMuxOut[1] = fifoOut[25][6][w-1];
              unloadMuxOut[2] = fifoOut[0][5][w-1];
              unloadMuxOut[3] = fifoOut[1][5][w-1];
              unloadMuxOut[4] = fifoOut[2][5][w-1];
              unloadMuxOut[5] = fifoOut[3][5][w-1];
              unloadMuxOut[6] = fifoOut[4][5][w-1];
              unloadMuxOut[7] = fifoOut[5][5][w-1];
              unloadMuxOut[8] = fifoOut[6][5][w-1];
              unloadMuxOut[9] = fifoOut[7][5][w-1];
              unloadMuxOut[10] = fifoOut[8][5][w-1];
              unloadMuxOut[11] = fifoOut[9][5][w-1];
              unloadMuxOut[12] = fifoOut[10][5][w-1];
              unloadMuxOut[13] = fifoOut[11][5][w-1];
              unloadMuxOut[14] = fifoOut[12][5][w-1];
              unloadMuxOut[15] = fifoOut[13][5][w-1];
              unloadMuxOut[16] = fifoOut[14][5][w-1];
              unloadMuxOut[17] = fifoOut[15][5][w-1];
              unloadMuxOut[18] = fifoOut[16][5][w-1];
              unloadMuxOut[19] = fifoOut[17][5][w-1];
              unloadMuxOut[20] = fifoOut[18][5][w-1];
              unloadMuxOut[21] = fifoOut[19][5][w-1];
              unloadMuxOut[22] = fifoOut[20][5][w-1];
              unloadMuxOut[23] = fifoOut[21][5][w-1];
              unloadMuxOut[24] = fifoOut[22][5][w-1];
              unloadMuxOut[25] = fifoOut[23][5][w-1];
              unloadMuxOut[26] = fifoOut[24][5][w-1];
              unloadMuxOut[27] = fifoOut[25][5][w-1];
              unloadMuxOut[28] = fifoOut[0][4][w-1];
              unloadMuxOut[29] = fifoOut[1][4][w-1];
              unloadMuxOut[30] = fifoOut[2][4][w-1];
              unloadMuxOut[31] = fifoOut[3][4][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[4][5][w-1];
              unloadMuxOut[1] = fifoOut[5][5][w-1];
              unloadMuxOut[2] = fifoOut[6][5][w-1];
              unloadMuxOut[3] = fifoOut[7][5][w-1];
              unloadMuxOut[4] = fifoOut[8][5][w-1];
              unloadMuxOut[5] = fifoOut[9][5][w-1];
              unloadMuxOut[6] = fifoOut[10][5][w-1];
              unloadMuxOut[7] = fifoOut[11][5][w-1];
              unloadMuxOut[8] = fifoOut[12][5][w-1];
              unloadMuxOut[9] = fifoOut[13][5][w-1];
              unloadMuxOut[10] = fifoOut[14][5][w-1];
              unloadMuxOut[11] = fifoOut[15][5][w-1];
              unloadMuxOut[12] = fifoOut[16][5][w-1];
              unloadMuxOut[13] = fifoOut[17][5][w-1];
              unloadMuxOut[14] = fifoOut[18][5][w-1];
              unloadMuxOut[15] = fifoOut[19][5][w-1];
              unloadMuxOut[16] = fifoOut[20][5][w-1];
              unloadMuxOut[17] = fifoOut[21][5][w-1];
              unloadMuxOut[18] = fifoOut[22][5][w-1];
              unloadMuxOut[19] = fifoOut[23][5][w-1];
              unloadMuxOut[20] = fifoOut[24][5][w-1];
              unloadMuxOut[21] = fifoOut[25][5][w-1];
              unloadMuxOut[22] = fifoOut[0][4][w-1];
              unloadMuxOut[23] = fifoOut[1][4][w-1];
              unloadMuxOut[24] = fifoOut[2][4][w-1];
              unloadMuxOut[25] = fifoOut[3][4][w-1];
              unloadMuxOut[26] = fifoOut[4][4][w-1];
              unloadMuxOut[27] = fifoOut[5][4][w-1];
              unloadMuxOut[28] = fifoOut[6][4][w-1];
              unloadMuxOut[29] = fifoOut[7][4][w-1];
              unloadMuxOut[30] = fifoOut[8][4][w-1];
              unloadMuxOut[31] = fifoOut[9][4][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[10][5][w-1];
              unloadMuxOut[1] = fifoOut[11][5][w-1];
              unloadMuxOut[2] = fifoOut[12][5][w-1];
              unloadMuxOut[3] = fifoOut[13][5][w-1];
              unloadMuxOut[4] = fifoOut[14][5][w-1];
              unloadMuxOut[5] = fifoOut[15][5][w-1];
              unloadMuxOut[6] = fifoOut[16][5][w-1];
              unloadMuxOut[7] = fifoOut[17][5][w-1];
              unloadMuxOut[8] = fifoOut[18][5][w-1];
              unloadMuxOut[9] = fifoOut[19][5][w-1];
              unloadMuxOut[10] = fifoOut[20][5][w-1];
              unloadMuxOut[11] = fifoOut[21][5][w-1];
              unloadMuxOut[12] = fifoOut[22][5][w-1];
              unloadMuxOut[13] = fifoOut[23][5][w-1];
              unloadMuxOut[14] = fifoOut[24][5][w-1];
              unloadMuxOut[15] = fifoOut[25][5][w-1];
              unloadMuxOut[16] = fifoOut[0][4][w-1];
              unloadMuxOut[17] = fifoOut[1][4][w-1];
              unloadMuxOut[18] = fifoOut[2][4][w-1];
              unloadMuxOut[19] = fifoOut[3][4][w-1];
              unloadMuxOut[20] = fifoOut[4][4][w-1];
              unloadMuxOut[21] = fifoOut[5][4][w-1];
              unloadMuxOut[22] = fifoOut[6][4][w-1];
              unloadMuxOut[23] = fifoOut[7][4][w-1];
              unloadMuxOut[24] = fifoOut[8][4][w-1];
              unloadMuxOut[25] = fifoOut[9][4][w-1];
              unloadMuxOut[26] = fifoOut[10][4][w-1];
              unloadMuxOut[27] = fifoOut[11][4][w-1];
              unloadMuxOut[28] = fifoOut[12][4][w-1];
              unloadMuxOut[29] = fifoOut[13][4][w-1];
              unloadMuxOut[30] = fifoOut[14][4][w-1];
              unloadMuxOut[31] = fifoOut[15][4][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[16][5][w-1];
              unloadMuxOut[1] = fifoOut[38][1][w-1];
              unloadMuxOut[2] = fifoOut[39][1][w-1];
              unloadMuxOut[3] = fifoOut[40][1][w-1];
              unloadMuxOut[4] = fifoOut[41][1][w-1];
              unloadMuxOut[5] = fifoOut[42][1][w-1];
              unloadMuxOut[6] = fifoOut[43][1][w-1];
              unloadMuxOut[7] = fifoOut[44][1][w-1];
              unloadMuxOut[8] = fifoOut[45][1][w-1];
              unloadMuxOut[9] = fifoOut[46][1][w-1];
              unloadMuxOut[10] = fifoOut[47][1][w-1];
              unloadMuxOut[11] = fifoOut[48][1][w-1];
              unloadMuxOut[12] = fifoOut[49][1][w-1];
              unloadMuxOut[13] = fifoOut[50][1][w-1];
              unloadMuxOut[14] = fifoOut[51][1][w-1];
              unloadMuxOut[15] = fifoOut[26][0][w-1];
              unloadMuxOut[16] = fifoOut[27][0][w-1];
              unloadMuxOut[17] = fifoOut[28][0][w-1];
              unloadMuxOut[18] = fifoOut[29][0][w-1];
              unloadMuxOut[19] = fifoOut[30][0][w-1];
              unloadMuxOut[20] = fifoOut[31][0][w-1];
              unloadMuxOut[21] = fifoOut[32][0][w-1];
              unloadMuxOut[22] = fifoOut[33][0][w-1];
              unloadMuxOut[23] = fifoOut[34][0][w-1];
              unloadMuxOut[24] = fifoOut[35][0][w-1];
              unloadMuxOut[25] = fifoOut[36][0][w-1];
              unloadMuxOut[26] = fifoOut[37][0][w-1];
              unloadMuxOut[27] = fifoOut[38][0][w-1];
              unloadMuxOut[28] = fifoOut[39][0][w-1];
              unloadMuxOut[29] = fifoOut[40][0][w-1];
              unloadMuxOut[30] = fifoOut[41][0][w-1];
              unloadMuxOut[31] = fifoOut[42][0][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[43][1][w-1];
              unloadMuxOut[1] = fifoOut[44][1][w-1];
              unloadMuxOut[2] = fifoOut[45][1][w-1];
              unloadMuxOut[3] = fifoOut[46][1][w-1];
              unloadMuxOut[4] = fifoOut[47][1][w-1];
              unloadMuxOut[5] = fifoOut[48][1][w-1];
              unloadMuxOut[6] = fifoOut[49][1][w-1];
              unloadMuxOut[7] = fifoOut[50][1][w-1];
              unloadMuxOut[8] = fifoOut[51][1][w-1];
              unloadMuxOut[9] = fifoOut[26][0][w-1];
              unloadMuxOut[10] = fifoOut[27][0][w-1];
              unloadMuxOut[11] = fifoOut[28][0][w-1];
              unloadMuxOut[12] = fifoOut[29][0][w-1];
              unloadMuxOut[13] = fifoOut[30][0][w-1];
              unloadMuxOut[14] = fifoOut[31][0][w-1];
              unloadMuxOut[15] = fifoOut[32][0][w-1];
              unloadMuxOut[16] = fifoOut[33][0][w-1];
              unloadMuxOut[17] = fifoOut[34][0][w-1];
              unloadMuxOut[18] = fifoOut[35][0][w-1];
              unloadMuxOut[19] = fifoOut[36][0][w-1];
              unloadMuxOut[20] = fifoOut[37][0][w-1];
              unloadMuxOut[21] = fifoOut[38][0][w-1];
              unloadMuxOut[22] = fifoOut[39][0][w-1];
              unloadMuxOut[23] = fifoOut[40][0][w-1];
              unloadMuxOut[24] = fifoOut[41][0][w-1];
              unloadMuxOut[25] = fifoOut[42][0][w-1];
              unloadMuxOut[26] = fifoOut[43][0][w-1];
              unloadMuxOut[27] = fifoOut[44][0][w-1];
              unloadMuxOut[28] = fifoOut[45][0][w-1];
              unloadMuxOut[29] = fifoOut[46][0][w-1];
              unloadMuxOut[30] = fifoOut[47][0][w-1];
              unloadMuxOut[31] = fifoOut[48][0][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[49][1][w-1];
              unloadMuxOut[1] = fifoOut[50][1][w-1];
              unloadMuxOut[2] = fifoOut[51][1][w-1];
              unloadMuxOut[3] = fifoOut[26][0][w-1];
              unloadMuxOut[4] = fifoOut[27][0][w-1];
              unloadMuxOut[5] = fifoOut[28][0][w-1];
              unloadMuxOut[6] = fifoOut[29][0][w-1];
              unloadMuxOut[7] = fifoOut[30][0][w-1];
              unloadMuxOut[8] = fifoOut[31][0][w-1];
              unloadMuxOut[9] = fifoOut[32][0][w-1];
              unloadMuxOut[10] = fifoOut[33][0][w-1];
              unloadMuxOut[11] = fifoOut[34][0][w-1];
              unloadMuxOut[12] = fifoOut[35][0][w-1];
              unloadMuxOut[13] = fifoOut[36][0][w-1];
              unloadMuxOut[14] = fifoOut[37][0][w-1];
              unloadMuxOut[15] = fifoOut[38][0][w-1];
              unloadMuxOut[16] = fifoOut[39][0][w-1];
              unloadMuxOut[17] = fifoOut[40][0][w-1];
              unloadMuxOut[18] = fifoOut[41][0][w-1];
              unloadMuxOut[19] = fifoOut[42][0][w-1];
              unloadMuxOut[20] = fifoOut[43][0][w-1];
              unloadMuxOut[21] = fifoOut[44][0][w-1];
              unloadMuxOut[22] = fifoOut[45][0][w-1];
              unloadMuxOut[23] = fifoOut[46][0][w-1];
              unloadMuxOut[24] = fifoOut[47][0][w-1];
              unloadMuxOut[25] = fifoOut[48][0][w-1];
              unloadMuxOut[26] = fifoOut[49][0][w-1];
              unloadMuxOut[27] = fifoOut[50][0][w-1];
              unloadMuxOut[28] = fifoOut[51][0][w-1];
              unloadMuxOut[29] = fifoOut[26][16][w-1];
              unloadMuxOut[30] = fifoOut[27][16][w-1];
              unloadMuxOut[31] = fifoOut[28][16][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[29][0][w-1];
              unloadMuxOut[1] = fifoOut[30][0][w-1];
              unloadMuxOut[2] = fifoOut[31][0][w-1];
              unloadMuxOut[3] = fifoOut[32][0][w-1];
              unloadMuxOut[4] = fifoOut[33][0][w-1];
              unloadMuxOut[5] = fifoOut[34][0][w-1];
              unloadMuxOut[6] = fifoOut[35][0][w-1];
              unloadMuxOut[7] = fifoOut[36][0][w-1];
              unloadMuxOut[8] = fifoOut[37][0][w-1];
              unloadMuxOut[9] = fifoOut[38][0][w-1];
              unloadMuxOut[10] = fifoOut[39][0][w-1];
              unloadMuxOut[11] = fifoOut[40][0][w-1];
              unloadMuxOut[12] = fifoOut[41][0][w-1];
              unloadMuxOut[13] = fifoOut[42][0][w-1];
              unloadMuxOut[14] = fifoOut[43][0][w-1];
              unloadMuxOut[15] = fifoOut[44][0][w-1];
              unloadMuxOut[16] = fifoOut[45][0][w-1];
              unloadMuxOut[17] = fifoOut[46][0][w-1];
              unloadMuxOut[18] = fifoOut[47][0][w-1];
              unloadMuxOut[19] = fifoOut[48][0][w-1];
              unloadMuxOut[20] = fifoOut[49][0][w-1];
              unloadMuxOut[21] = fifoOut[50][0][w-1];
              unloadMuxOut[22] = fifoOut[51][0][w-1];
              unloadMuxOut[23] = fifoOut[26][16][w-1];
              unloadMuxOut[24] = fifoOut[27][16][w-1];
              unloadMuxOut[25] = fifoOut[28][16][w-1];
              unloadMuxOut[26] = fifoOut[29][16][w-1];
              unloadMuxOut[27] = fifoOut[30][16][w-1];
              unloadMuxOut[28] = fifoOut[31][16][w-1];
              unloadMuxOut[29] = fifoOut[32][16][w-1];
              unloadMuxOut[30] = fifoOut[33][16][w-1];
              unloadMuxOut[31] = fifoOut[34][16][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[35][0][w-1];
              unloadMuxOut[1] = fifoOut[36][0][w-1];
              unloadMuxOut[2] = fifoOut[37][0][w-1];
              unloadMuxOut[3] = fifoOut[38][0][w-1];
              unloadMuxOut[4] = fifoOut[39][0][w-1];
              unloadMuxOut[5] = fifoOut[40][0][w-1];
              unloadMuxOut[6] = fifoOut[41][0][w-1];
              unloadMuxOut[7] = fifoOut[42][0][w-1];
              unloadMuxOut[8] = fifoOut[43][0][w-1];
              unloadMuxOut[9] = fifoOut[44][0][w-1];
              unloadMuxOut[10] = fifoOut[45][0][w-1];
              unloadMuxOut[11] = fifoOut[46][0][w-1];
              unloadMuxOut[12] = fifoOut[47][0][w-1];
              unloadMuxOut[13] = fifoOut[48][0][w-1];
              unloadMuxOut[14] = fifoOut[49][0][w-1];
              unloadMuxOut[15] = fifoOut[50][0][w-1];
              unloadMuxOut[16] = fifoOut[51][0][w-1];
              unloadMuxOut[17] = fifoOut[26][16][w-1];
              unloadMuxOut[18] = fifoOut[27][16][w-1];
              unloadMuxOut[19] = fifoOut[28][16][w-1];
              unloadMuxOut[20] = fifoOut[29][16][w-1];
              unloadMuxOut[21] = fifoOut[30][16][w-1];
              unloadMuxOut[22] = fifoOut[31][16][w-1];
              unloadMuxOut[23] = fifoOut[32][16][w-1];
              unloadMuxOut[24] = fifoOut[33][16][w-1];
              unloadMuxOut[25] = fifoOut[34][16][w-1];
              unloadMuxOut[26] = fifoOut[35][16][w-1];
              unloadMuxOut[27] = fifoOut[36][16][w-1];
              unloadMuxOut[28] = fifoOut[37][16][w-1];
              unloadMuxOut[29] = fifoOut[38][16][w-1];
              unloadMuxOut[30] = fifoOut[39][16][w-1];
              unloadMuxOut[31] = fifoOut[40][16][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[3][6][w-1];
              unloadMuxOut[1] = fifoOut[4][6][w-1];
              unloadMuxOut[2] = fifoOut[5][6][w-1];
              unloadMuxOut[3] = fifoOut[6][6][w-1];
              unloadMuxOut[4] = fifoOut[7][6][w-1];
              unloadMuxOut[5] = fifoOut[8][6][w-1];
              unloadMuxOut[6] = fifoOut[9][6][w-1];
              unloadMuxOut[7] = fifoOut[10][6][w-1];
              unloadMuxOut[8] = fifoOut[11][6][w-1];
              unloadMuxOut[9] = fifoOut[12][6][w-1];
              unloadMuxOut[10] = fifoOut[13][6][w-1];
              unloadMuxOut[11] = fifoOut[26][16][w-1];
              unloadMuxOut[12] = fifoOut[27][16][w-1];
              unloadMuxOut[13] = fifoOut[28][16][w-1];
              unloadMuxOut[14] = fifoOut[29][16][w-1];
              unloadMuxOut[15] = fifoOut[30][16][w-1];
              unloadMuxOut[16] = fifoOut[31][16][w-1];
              unloadMuxOut[17] = fifoOut[32][16][w-1];
              unloadMuxOut[18] = fifoOut[33][16][w-1];
              unloadMuxOut[19] = fifoOut[34][16][w-1];
              unloadMuxOut[20] = fifoOut[35][16][w-1];
              unloadMuxOut[21] = fifoOut[36][16][w-1];
              unloadMuxOut[22] = fifoOut[37][16][w-1];
              unloadMuxOut[23] = fifoOut[38][16][w-1];
              unloadMuxOut[24] = fifoOut[39][16][w-1];
              unloadMuxOut[25] = fifoOut[40][16][w-1];
              unloadMuxOut[26] = fifoOut[41][16][w-1];
              unloadMuxOut[27] = fifoOut[42][16][w-1];
              unloadMuxOut[28] = fifoOut[43][16][w-1];
              unloadMuxOut[29] = fifoOut[44][16][w-1];
              unloadMuxOut[30] = fifoOut[45][16][w-1];
              unloadMuxOut[31] = fifoOut[46][16][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[9][6][w-1];
              unloadMuxOut[1] = fifoOut[10][6][w-1];
              unloadMuxOut[2] = fifoOut[11][6][w-1];
              unloadMuxOut[3] = fifoOut[12][6][w-1];
              unloadMuxOut[4] = fifoOut[13][6][w-1];
              unloadMuxOut[5] = fifoOut[26][16][w-1];
              unloadMuxOut[6] = fifoOut[27][16][w-1];
              unloadMuxOut[7] = fifoOut[28][16][w-1];
              unloadMuxOut[8] = fifoOut[29][16][w-1];
              unloadMuxOut[9] = fifoOut[30][16][w-1];
              unloadMuxOut[10] = fifoOut[31][16][w-1];
              unloadMuxOut[11] = fifoOut[32][16][w-1];
              unloadMuxOut[12] = fifoOut[33][16][w-1];
              unloadMuxOut[13] = fifoOut[34][16][w-1];
              unloadMuxOut[14] = fifoOut[35][16][w-1];
              unloadMuxOut[15] = fifoOut[36][16][w-1];
              unloadMuxOut[16] = fifoOut[37][16][w-1];
              unloadMuxOut[17] = fifoOut[38][16][w-1];
              unloadMuxOut[18] = fifoOut[39][16][w-1];
              unloadMuxOut[19] = fifoOut[40][16][w-1];
              unloadMuxOut[20] = fifoOut[41][16][w-1];
              unloadMuxOut[21] = fifoOut[42][16][w-1];
              unloadMuxOut[22] = fifoOut[43][16][w-1];
              unloadMuxOut[23] = fifoOut[44][16][w-1];
              unloadMuxOut[24] = fifoOut[45][16][w-1];
              unloadMuxOut[25] = fifoOut[46][16][w-1];
              unloadMuxOut[26] = fifoOut[47][16][w-1];
              unloadMuxOut[27] = fifoOut[48][16][w-1];
              unloadMuxOut[28] = fifoOut[49][16][w-1];
              unloadMuxOut[29] = fifoOut[50][16][w-1];
              unloadMuxOut[30] = fifoOut[51][16][w-1];
              unloadMuxOut[31] = fifoOut[26][15][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[27][16][w-1];
              unloadMuxOut[1] = fifoOut[28][16][w-1];
              unloadMuxOut[2] = fifoOut[29][16][w-1];
              unloadMuxOut[3] = fifoOut[30][16][w-1];
              unloadMuxOut[4] = fifoOut[31][16][w-1];
              unloadMuxOut[5] = fifoOut[32][16][w-1];
              unloadMuxOut[6] = fifoOut[33][16][w-1];
              unloadMuxOut[7] = fifoOut[34][16][w-1];
              unloadMuxOut[8] = fifoOut[35][16][w-1];
              unloadMuxOut[9] = fifoOut[36][16][w-1];
              unloadMuxOut[10] = fifoOut[37][16][w-1];
              unloadMuxOut[11] = fifoOut[38][16][w-1];
              unloadMuxOut[12] = fifoOut[39][16][w-1];
              unloadMuxOut[13] = fifoOut[40][16][w-1];
              unloadMuxOut[14] = fifoOut[41][16][w-1];
              unloadMuxOut[15] = fifoOut[42][16][w-1];
              unloadMuxOut[16] = fifoOut[43][16][w-1];
              unloadMuxOut[17] = fifoOut[44][16][w-1];
              unloadMuxOut[18] = fifoOut[45][16][w-1];
              unloadMuxOut[19] = fifoOut[46][16][w-1];
              unloadMuxOut[20] = fifoOut[47][16][w-1];
              unloadMuxOut[21] = fifoOut[48][16][w-1];
              unloadMuxOut[22] = fifoOut[49][16][w-1];
              unloadMuxOut[23] = fifoOut[50][16][w-1];
              unloadMuxOut[24] = fifoOut[51][16][w-1];
              unloadMuxOut[25] = fifoOut[26][15][w-1];
              unloadMuxOut[26] = fifoOut[27][15][w-1];
              unloadMuxOut[27] = fifoOut[28][15][w-1];
              unloadMuxOut[28] = fifoOut[29][15][w-1];
              unloadMuxOut[29] = fifoOut[30][15][w-1];
              unloadMuxOut[30] = fifoOut[31][15][w-1];
              unloadMuxOut[31] = fifoOut[32][15][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[33][16][w-1];
              unloadMuxOut[1] = fifoOut[34][16][w-1];
              unloadMuxOut[2] = fifoOut[35][16][w-1];
              unloadMuxOut[3] = fifoOut[36][16][w-1];
              unloadMuxOut[4] = fifoOut[37][16][w-1];
              unloadMuxOut[5] = fifoOut[38][16][w-1];
              unloadMuxOut[6] = fifoOut[39][16][w-1];
              unloadMuxOut[7] = fifoOut[40][16][w-1];
              unloadMuxOut[8] = fifoOut[41][16][w-1];
              unloadMuxOut[9] = fifoOut[42][16][w-1];
              unloadMuxOut[10] = fifoOut[43][16][w-1];
              unloadMuxOut[11] = fifoOut[44][16][w-1];
              unloadMuxOut[12] = fifoOut[45][16][w-1];
              unloadMuxOut[13] = fifoOut[46][16][w-1];
              unloadMuxOut[14] = fifoOut[47][16][w-1];
              unloadMuxOut[15] = fifoOut[48][16][w-1];
              unloadMuxOut[16] = fifoOut[49][16][w-1];
              unloadMuxOut[17] = fifoOut[50][16][w-1];
              unloadMuxOut[18] = fifoOut[51][16][w-1];
              unloadMuxOut[19] = fifoOut[26][15][w-1];
              unloadMuxOut[20] = fifoOut[27][15][w-1];
              unloadMuxOut[21] = fifoOut[28][15][w-1];
              unloadMuxOut[22] = fifoOut[29][15][w-1];
              unloadMuxOut[23] = fifoOut[30][15][w-1];
              unloadMuxOut[24] = fifoOut[31][15][w-1];
              unloadMuxOut[25] = fifoOut[32][15][w-1];
              unloadMuxOut[26] = fifoOut[33][15][w-1];
              unloadMuxOut[27] = fifoOut[34][15][w-1];
              unloadMuxOut[28] = fifoOut[35][15][w-1];
              unloadMuxOut[29] = fifoOut[36][15][w-1];
              unloadMuxOut[30] = fifoOut[37][15][w-1];
              unloadMuxOut[31] = fifoOut[38][15][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[39][16][w-1];
              unloadMuxOut[1] = fifoOut[40][16][w-1];
              unloadMuxOut[2] = fifoOut[41][16][w-1];
              unloadMuxOut[3] = fifoOut[42][16][w-1];
              unloadMuxOut[4] = fifoOut[43][16][w-1];
              unloadMuxOut[5] = fifoOut[44][16][w-1];
              unloadMuxOut[6] = fifoOut[45][16][w-1];
              unloadMuxOut[7] = fifoOut[46][16][w-1];
              unloadMuxOut[8] = fifoOut[47][16][w-1];
              unloadMuxOut[9] = fifoOut[48][16][w-1];
              unloadMuxOut[10] = fifoOut[49][16][w-1];
              unloadMuxOut[11] = fifoOut[50][16][w-1];
              unloadMuxOut[12] = fifoOut[51][16][w-1];
              unloadMuxOut[13] = fifoOut[26][15][w-1];
              unloadMuxOut[14] = fifoOut[27][15][w-1];
              unloadMuxOut[15] = fifoOut[28][15][w-1];
              unloadMuxOut[16] = fifoOut[29][15][w-1];
              unloadMuxOut[17] = fifoOut[30][15][w-1];
              unloadMuxOut[18] = fifoOut[31][15][w-1];
              unloadMuxOut[19] = fifoOut[32][15][w-1];
              unloadMuxOut[20] = fifoOut[33][15][w-1];
              unloadMuxOut[21] = fifoOut[34][15][w-1];
              unloadMuxOut[22] = fifoOut[35][15][w-1];
              unloadMuxOut[23] = fifoOut[36][15][w-1];
              unloadMuxOut[24] = fifoOut[37][15][w-1];
              unloadMuxOut[25] = fifoOut[38][15][w-1];
              unloadMuxOut[26] = fifoOut[39][15][w-1];
              unloadMuxOut[27] = fifoOut[40][15][w-1];
              unloadMuxOut[28] = fifoOut[41][15][w-1];
              unloadMuxOut[29] = fifoOut[42][15][w-1];
              unloadMuxOut[30] = fifoOut[43][15][w-1];
              unloadMuxOut[31] = fifoOut[44][15][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[45][16][w-1];
              unloadMuxOut[1] = fifoOut[46][16][w-1];
              unloadMuxOut[2] = fifoOut[47][16][w-1];
              unloadMuxOut[3] = fifoOut[48][16][w-1];
              unloadMuxOut[4] = fifoOut[49][16][w-1];
              unloadMuxOut[5] = fifoOut[50][16][w-1];
              unloadMuxOut[6] = fifoOut[51][16][w-1];
              unloadMuxOut[7] = fifoOut[26][15][w-1];
              unloadMuxOut[8] = fifoOut[27][15][w-1];
              unloadMuxOut[9] = fifoOut[28][15][w-1];
              unloadMuxOut[10] = fifoOut[29][15][w-1];
              unloadMuxOut[11] = fifoOut[30][15][w-1];
              unloadMuxOut[12] = fifoOut[31][15][w-1];
              unloadMuxOut[13] = fifoOut[32][15][w-1];
              unloadMuxOut[14] = fifoOut[33][15][w-1];
              unloadMuxOut[15] = fifoOut[34][15][w-1];
              unloadMuxOut[16] = fifoOut[35][15][w-1];
              unloadMuxOut[17] = fifoOut[36][15][w-1];
              unloadMuxOut[18] = fifoOut[37][15][w-1];
              unloadMuxOut[19] = fifoOut[38][15][w-1];
              unloadMuxOut[20] = fifoOut[39][15][w-1];
              unloadMuxOut[21] = fifoOut[40][15][w-1];
              unloadMuxOut[22] = fifoOut[41][15][w-1];
              unloadMuxOut[23] = fifoOut[42][15][w-1];
              unloadMuxOut[24] = fifoOut[5][4][w-1];
              unloadMuxOut[25] = fifoOut[6][4][w-1];
              unloadMuxOut[26] = fifoOut[7][4][w-1];
              unloadMuxOut[27] = fifoOut[8][4][w-1];
              unloadMuxOut[28] = fifoOut[9][4][w-1];
              unloadMuxOut[29] = fifoOut[10][4][w-1];
              unloadMuxOut[30] = fifoOut[11][4][w-1];
              unloadMuxOut[31] = fifoOut[12][4][w-1];
       end
       16: begin
              unloadMuxOut[0] = fifoOut[13][5][w-1];
              unloadMuxOut[1] = fifoOut[14][5][w-1];
              unloadMuxOut[2] = fifoOut[15][5][w-1];
              unloadMuxOut[3] = fifoOut[16][5][w-1];
              unloadMuxOut[4] = fifoOut[17][5][w-1];
              unloadMuxOut[5] = fifoOut[18][5][w-1];
              unloadMuxOut[6] = fifoOut[19][5][w-1];
              unloadMuxOut[7] = fifoOut[20][5][w-1];
              unloadMuxOut[8] = fifoOut[21][5][w-1];
              unloadMuxOut[9] = fifoOut[22][5][w-1];
              unloadMuxOut[10] = fifoOut[23][5][w-1];
              unloadMuxOut[11] = fifoOut[24][5][w-1];
              unloadMuxOut[12] = fifoOut[25][5][w-1];
              unloadMuxOut[13] = fifoOut[0][4][w-1];
              unloadMuxOut[14] = fifoOut[1][4][w-1];
              unloadMuxOut[15] = fifoOut[2][4][w-1];
              unloadMuxOut[16] = fifoOut[3][4][w-1];
              unloadMuxOut[17] = fifoOut[4][4][w-1];
              unloadMuxOut[18] = fifoOut[5][4][w-1];
              unloadMuxOut[19] = fifoOut[6][4][w-1];
              unloadMuxOut[20] = fifoOut[7][4][w-1];
              unloadMuxOut[21] = fifoOut[8][4][w-1];
              unloadMuxOut[22] = fifoOut[9][4][w-1];
              unloadMuxOut[23] = fifoOut[10][4][w-1];
              unloadMuxOut[24] = fifoOut[11][4][w-1];
              unloadMuxOut[25] = fifoOut[12][4][w-1];
              unloadMuxOut[26] = fifoOut[13][4][w-1];
              unloadMuxOut[27] = fifoOut[14][4][w-1];
              unloadMuxOut[28] = fifoOut[15][4][w-1];
              unloadMuxOut[29] = fifoOut[16][4][w-1];
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0; 
             end
       end
    endcase //unload case end
    case(iteration_0_indicator)
       0: begin
         case(rd_address_case)
         0: begin
              muxOutConnector[0] = fifoOut[3][4];
              muxOutConnector[1] = fifoOut[4][4];
              muxOutConnector[2] = fifoOut[5][4];
              muxOutConnector[3] = fifoOut[6][4];
              muxOutConnector[4] = fifoOut[7][4];
              muxOutConnector[5] = fifoOut[8][4];
              muxOutConnector[6] = fifoOut[9][4];
              muxOutConnector[7] = fifoOut[10][4];
              muxOutConnector[8] = fifoOut[11][4];
              muxOutConnector[9] = fifoOut[12][4];
              muxOutConnector[10] = fifoOut[13][4];
              muxOutConnector[11] = fifoOut[14][4];
              muxOutConnector[12] = fifoOut[15][4];
              muxOutConnector[13] = fifoOut[16][4];
              muxOutConnector[14] = fifoOut[17][4];
              muxOutConnector[15] = fifoOut[18][4];
              muxOutConnector[16] = fifoOut[19][4];
              muxOutConnector[17] = fifoOut[20][4];
              muxOutConnector[18] = fifoOut[21][4];
              muxOutConnector[19] = fifoOut[22][4];
              muxOutConnector[20] = fifoOut[23][4];
              muxOutConnector[21] = fifoOut[24][4];
              muxOutConnector[22] = fifoOut[25][4];
              muxOutConnector[23] = fifoOut[0][3];
              muxOutConnector[24] = fifoOut[1][3];
              muxOutConnector[25] = fifoOut[2][3];
              muxOutConnector[26] = fifoOut[43][9];
              muxOutConnector[27] = fifoOut[44][9];
              muxOutConnector[28] = fifoOut[45][9];
              muxOutConnector[29] = fifoOut[46][9];
              muxOutConnector[30] = fifoOut[47][9];
              muxOutConnector[31] = fifoOut[48][9];
              muxOutConnector[32] = fifoOut[49][9];
              muxOutConnector[33] = fifoOut[50][9];
              muxOutConnector[34] = fifoOut[51][9];
              muxOutConnector[35] = fifoOut[26][8];
              muxOutConnector[36] = fifoOut[27][8];
              muxOutConnector[37] = fifoOut[28][8];
              muxOutConnector[38] = fifoOut[29][8];
              muxOutConnector[39] = fifoOut[30][8];
              muxOutConnector[40] = fifoOut[31][8];
              muxOutConnector[41] = fifoOut[32][8];
              muxOutConnector[42] = fifoOut[33][8];
              muxOutConnector[43] = fifoOut[34][8];
              muxOutConnector[44] = fifoOut[35][8];
              muxOutConnector[45] = fifoOut[36][8];
              muxOutConnector[46] = fifoOut[37][8];
              muxOutConnector[47] = fifoOut[38][8];
              muxOutConnector[48] = fifoOut[39][8];
              muxOutConnector[49] = fifoOut[40][8];
              muxOutConnector[50] = fifoOut[41][8];
              muxOutConnector[51] = fifoOut[42][8];
         end
         1: begin
              muxOutConnector[0] = fifoOut[3][4];
              muxOutConnector[1] = fifoOut[4][4];
              muxOutConnector[2] = fifoOut[5][4];
              muxOutConnector[3] = fifoOut[6][4];
              muxOutConnector[4] = fifoOut[7][4];
              muxOutConnector[5] = fifoOut[8][4];
              muxOutConnector[6] = fifoOut[9][4];
              muxOutConnector[7] = fifoOut[10][4];
              muxOutConnector[8] = fifoOut[11][4];
              muxOutConnector[9] = fifoOut[12][4];
              muxOutConnector[10] = fifoOut[13][4];
              muxOutConnector[11] = fifoOut[14][4];
              muxOutConnector[12] = fifoOut[15][4];
              muxOutConnector[13] = fifoOut[16][4];
              muxOutConnector[14] = fifoOut[17][4];
              muxOutConnector[15] = fifoOut[18][4];
              muxOutConnector[16] = fifoOut[19][4];
              muxOutConnector[17] = fifoOut[20][4];
              muxOutConnector[18] = fifoOut[21][4];
              muxOutConnector[19] = fifoOut[22][4];
              muxOutConnector[20] = fifoOut[23][4];
              muxOutConnector[21] = fifoOut[24][4];
              muxOutConnector[22] = fifoOut[25][4];
              muxOutConnector[23] = fifoOut[0][3];
              muxOutConnector[24] = fifoOut[1][3];
              muxOutConnector[25] = fifoOut[2][3];
              muxOutConnector[26] = fifoOut[43][9];
              muxOutConnector[27] = fifoOut[44][9];
              muxOutConnector[28] = fifoOut[45][9];
              muxOutConnector[29] = fifoOut[46][9];
              muxOutConnector[30] = fifoOut[47][9];
              muxOutConnector[31] = fifoOut[48][9];
              muxOutConnector[32] = fifoOut[49][9];
              muxOutConnector[33] = fifoOut[50][9];
              muxOutConnector[34] = fifoOut[51][9];
              muxOutConnector[35] = fifoOut[26][8];
              muxOutConnector[36] = fifoOut[27][8];
              muxOutConnector[37] = fifoOut[28][8];
              muxOutConnector[38] = fifoOut[29][8];
              muxOutConnector[39] = fifoOut[30][8];
              muxOutConnector[40] = fifoOut[31][8];
              muxOutConnector[41] = fifoOut[32][8];
              muxOutConnector[42] = fifoOut[33][8];
              muxOutConnector[43] = fifoOut[34][8];
              muxOutConnector[44] = fifoOut[35][8];
              muxOutConnector[45] = fifoOut[36][8];
              muxOutConnector[46] = fifoOut[37][8];
              muxOutConnector[47] = fifoOut[0][14];
              muxOutConnector[48] = fifoOut[1][14];
              muxOutConnector[49] = fifoOut[2][14];
              muxOutConnector[50] = fifoOut[3][14];
              muxOutConnector[51] = fifoOut[4][14];
         end
         2: begin
              muxOutConnector[0] = fifoOut[3][4];
              muxOutConnector[1] = fifoOut[4][4];
              muxOutConnector[2] = fifoOut[5][4];
              muxOutConnector[3] = fifoOut[6][4];
              muxOutConnector[4] = fifoOut[7][4];
              muxOutConnector[5] = fifoOut[8][4];
              muxOutConnector[6] = fifoOut[9][4];
              muxOutConnector[7] = fifoOut[10][4];
              muxOutConnector[8] = fifoOut[11][4];
              muxOutConnector[9] = fifoOut[12][4];
              muxOutConnector[10] = fifoOut[13][4];
              muxOutConnector[11] = fifoOut[14][4];
              muxOutConnector[12] = fifoOut[15][4];
              muxOutConnector[13] = fifoOut[16][4];
              muxOutConnector[14] = fifoOut[17][4];
              muxOutConnector[15] = fifoOut[18][4];
              muxOutConnector[16] = fifoOut[19][4];
              muxOutConnector[17] = fifoOut[20][4];
              muxOutConnector[18] = fifoOut[21][4];
              muxOutConnector[19] = fifoOut[22][4];
              muxOutConnector[20] = fifoOut[23][4];
              muxOutConnector[21] = fifoOut[24][4];
              muxOutConnector[22] = fifoOut[25][4];
              muxOutConnector[23] = fifoOut[0][3];
              muxOutConnector[24] = fifoOut[1][3];
              muxOutConnector[25] = fifoOut[2][3];
              muxOutConnector[26] = fifoOut[5][15];
              muxOutConnector[27] = fifoOut[6][15];
              muxOutConnector[28] = fifoOut[7][15];
              muxOutConnector[29] = fifoOut[8][15];
              muxOutConnector[30] = fifoOut[9][15];
              muxOutConnector[31] = fifoOut[10][15];
              muxOutConnector[32] = fifoOut[11][15];
              muxOutConnector[33] = fifoOut[12][15];
              muxOutConnector[34] = fifoOut[13][15];
              muxOutConnector[35] = fifoOut[14][15];
              muxOutConnector[36] = fifoOut[15][15];
              muxOutConnector[37] = fifoOut[16][15];
              muxOutConnector[38] = fifoOut[17][15];
              muxOutConnector[39] = fifoOut[18][15];
              muxOutConnector[40] = fifoOut[19][15];
              muxOutConnector[41] = fifoOut[20][15];
              muxOutConnector[42] = fifoOut[21][15];
              muxOutConnector[43] = fifoOut[22][15];
              muxOutConnector[44] = fifoOut[23][15];
              muxOutConnector[45] = fifoOut[24][15];
              muxOutConnector[46] = fifoOut[25][15];
              muxOutConnector[47] = fifoOut[0][14];
              muxOutConnector[48] = fifoOut[1][14];
              muxOutConnector[49] = fifoOut[2][14];
              muxOutConnector[50] = fifoOut[3][14];
              muxOutConnector[51] = fifoOut[4][14];
         end
         3: begin
              muxOutConnector[0] = fifoOut[3][4];
              muxOutConnector[1] = fifoOut[4][4];
              muxOutConnector[2] = fifoOut[5][4];
              muxOutConnector[3] = fifoOut[6][4];
              muxOutConnector[4] = fifoOut[7][4];
              muxOutConnector[5] = fifoOut[8][4];
              muxOutConnector[6] = fifoOut[9][4];
              muxOutConnector[7] = fifoOut[10][4];
              muxOutConnector[8] = fifoOut[11][4];
              muxOutConnector[9] = fifoOut[12][4];
              muxOutConnector[10] = fifoOut[13][4];
              muxOutConnector[11] = fifoOut[14][4];
              muxOutConnector[12] = fifoOut[15][4];
              muxOutConnector[13] = fifoOut[16][4];
              muxOutConnector[14] = fifoOut[17][4];
              muxOutConnector[15] = fifoOut[18][4];
              muxOutConnector[16] = fifoOut[19][4];
              muxOutConnector[17] = fifoOut[20][4];
              muxOutConnector[18] = fifoOut[21][4];
              muxOutConnector[19] = fifoOut[22][4];
              muxOutConnector[20] = fifoOut[23][4];
              muxOutConnector[21] = fifoOut[24][4];
              muxOutConnector[22] = fifoOut[25][4];
              muxOutConnector[23] = fifoOut[0][3];
              muxOutConnector[24] = fifoOut[1][3];
              muxOutConnector[25] = fifoOut[2][3];
              muxOutConnector[26] = fifoOut[5][15];
              muxOutConnector[27] = fifoOut[6][15];
              muxOutConnector[28] = fifoOut[7][15];
              muxOutConnector[29] = fifoOut[8][15];
              muxOutConnector[30] = fifoOut[9][15];
              muxOutConnector[31] = fifoOut[10][15];
              muxOutConnector[32] = fifoOut[11][15];
              muxOutConnector[33] = fifoOut[12][15];
              muxOutConnector[34] = fifoOut[13][15];
              muxOutConnector[35] = fifoOut[14][15];
              muxOutConnector[36] = fifoOut[15][15];
              muxOutConnector[37] = fifoOut[16][15];
              muxOutConnector[38] = fifoOut[17][15];
              muxOutConnector[39] = fifoOut[18][15];
              muxOutConnector[40] = fifoOut[19][15];
              muxOutConnector[41] = fifoOut[20][15];
              muxOutConnector[42] = fifoOut[21][15];
              muxOutConnector[43] = fifoOut[22][15];
              muxOutConnector[44] = fifoOut[23][15];
              muxOutConnector[45] = fifoOut[24][15];
              muxOutConnector[46] = fifoOut[25][15];
              muxOutConnector[47] = fifoOut[0][14];
              muxOutConnector[48] = fifoOut[1][14];
              muxOutConnector[49] = fifoOut[2][14];
              muxOutConnector[50] = fifoOut[3][14];
              muxOutConnector[51] = fifoOut[4][14];
         end
         4: begin
              muxOutConnector[0] = fifoOut[3][4];
              muxOutConnector[1] = fifoOut[4][4];
              muxOutConnector[2] = fifoOut[5][4];
              muxOutConnector[3] = fifoOut[6][4];
              muxOutConnector[4] = fifoOut[7][4];
              muxOutConnector[5] = fifoOut[8][4];
              muxOutConnector[6] = fifoOut[9][4];
              muxOutConnector[7] = fifoOut[10][4];
              muxOutConnector[8] = fifoOut[11][4];
              muxOutConnector[9] = fifoOut[12][4];
              muxOutConnector[10] = fifoOut[13][4];
              muxOutConnector[11] = fifoOut[14][4];
              muxOutConnector[12] = fifoOut[15][4];
              muxOutConnector[13] = fifoOut[16][4];
              muxOutConnector[14] = fifoOut[38][0];
              muxOutConnector[15] = fifoOut[39][0];
              muxOutConnector[16] = fifoOut[40][0];
              muxOutConnector[17] = fifoOut[41][0];
              muxOutConnector[18] = fifoOut[42][0];
              muxOutConnector[19] = fifoOut[43][0];
              muxOutConnector[20] = fifoOut[44][0];
              muxOutConnector[21] = fifoOut[45][0];
              muxOutConnector[22] = fifoOut[46][0];
              muxOutConnector[23] = fifoOut[47][0];
              muxOutConnector[24] = fifoOut[48][0];
              muxOutConnector[25] = fifoOut[49][0];
              muxOutConnector[26] = fifoOut[5][15];
              muxOutConnector[27] = fifoOut[6][15];
              muxOutConnector[28] = fifoOut[7][15];
              muxOutConnector[29] = fifoOut[8][15];
              muxOutConnector[30] = fifoOut[9][15];
              muxOutConnector[31] = fifoOut[10][15];
              muxOutConnector[32] = fifoOut[11][15];
              muxOutConnector[33] = fifoOut[12][15];
              muxOutConnector[34] = fifoOut[13][15];
              muxOutConnector[35] = fifoOut[14][15];
              muxOutConnector[36] = fifoOut[15][15];
              muxOutConnector[37] = fifoOut[16][15];
              muxOutConnector[38] = fifoOut[17][15];
              muxOutConnector[39] = fifoOut[18][15];
              muxOutConnector[40] = fifoOut[19][15];
              muxOutConnector[41] = fifoOut[20][15];
              muxOutConnector[42] = fifoOut[21][15];
              muxOutConnector[43] = fifoOut[22][15];
              muxOutConnector[44] = fifoOut[23][15];
              muxOutConnector[45] = fifoOut[24][15];
              muxOutConnector[46] = fifoOut[25][15];
              muxOutConnector[47] = fifoOut[0][14];
              muxOutConnector[48] = fifoOut[1][14];
              muxOutConnector[49] = fifoOut[2][14];
              muxOutConnector[50] = fifoOut[3][14];
              muxOutConnector[51] = fifoOut[4][14];
         end
         5: begin
              muxOutConnector[0] = fifoOut[50][1];
              muxOutConnector[1] = fifoOut[51][1];
              muxOutConnector[2] = fifoOut[26][0];
              muxOutConnector[3] = fifoOut[27][0];
              muxOutConnector[4] = fifoOut[28][0];
              muxOutConnector[5] = fifoOut[29][0];
              muxOutConnector[6] = fifoOut[30][0];
              muxOutConnector[7] = fifoOut[31][0];
              muxOutConnector[8] = fifoOut[32][0];
              muxOutConnector[9] = fifoOut[33][0];
              muxOutConnector[10] = fifoOut[34][0];
              muxOutConnector[11] = fifoOut[35][0];
              muxOutConnector[12] = fifoOut[36][0];
              muxOutConnector[13] = fifoOut[37][0];
              muxOutConnector[14] = fifoOut[38][0];
              muxOutConnector[15] = fifoOut[39][0];
              muxOutConnector[16] = fifoOut[40][0];
              muxOutConnector[17] = fifoOut[41][0];
              muxOutConnector[18] = fifoOut[42][0];
              muxOutConnector[19] = fifoOut[43][0];
              muxOutConnector[20] = fifoOut[44][0];
              muxOutConnector[21] = fifoOut[45][0];
              muxOutConnector[22] = fifoOut[46][0];
              muxOutConnector[23] = fifoOut[47][0];
              muxOutConnector[24] = fifoOut[48][0];
              muxOutConnector[25] = fifoOut[49][0];
              muxOutConnector[26] = fifoOut[5][15];
              muxOutConnector[27] = fifoOut[6][15];
              muxOutConnector[28] = fifoOut[7][15];
              muxOutConnector[29] = fifoOut[8][15];
              muxOutConnector[30] = fifoOut[9][15];
              muxOutConnector[31] = fifoOut[10][15];
              muxOutConnector[32] = fifoOut[11][15];
              muxOutConnector[33] = fifoOut[12][15];
              muxOutConnector[34] = fifoOut[13][15];
              muxOutConnector[35] = fifoOut[14][15];
              muxOutConnector[36] = fifoOut[15][15];
              muxOutConnector[37] = fifoOut[16][15];
              muxOutConnector[38] = fifoOut[17][15];
              muxOutConnector[39] = fifoOut[18][15];
              muxOutConnector[40] = fifoOut[19][15];
              muxOutConnector[41] = fifoOut[20][15];
              muxOutConnector[42] = fifoOut[21][15];
              muxOutConnector[43] = fifoOut[22][15];
              muxOutConnector[44] = fifoOut[23][15];
              muxOutConnector[45] = fifoOut[24][15];
              muxOutConnector[46] = fifoOut[25][15];
              muxOutConnector[47] = fifoOut[0][14];
              muxOutConnector[48] = fifoOut[1][14];
              muxOutConnector[49] = fifoOut[2][14];
              muxOutConnector[50] = fifoOut[3][14];
              muxOutConnector[51] = fifoOut[4][14];
         end
         6: begin
              muxOutConnector[0] = fifoOut[50][1];
              muxOutConnector[1] = fifoOut[51][1];
              muxOutConnector[2] = fifoOut[26][0];
              muxOutConnector[3] = fifoOut[27][0];
              muxOutConnector[4] = fifoOut[28][0];
              muxOutConnector[5] = fifoOut[29][0];
              muxOutConnector[6] = fifoOut[30][0];
              muxOutConnector[7] = fifoOut[31][0];
              muxOutConnector[8] = fifoOut[32][0];
              muxOutConnector[9] = fifoOut[33][0];
              muxOutConnector[10] = fifoOut[34][0];
              muxOutConnector[11] = fifoOut[35][0];
              muxOutConnector[12] = fifoOut[36][0];
              muxOutConnector[13] = fifoOut[37][0];
              muxOutConnector[14] = fifoOut[38][0];
              muxOutConnector[15] = fifoOut[39][0];
              muxOutConnector[16] = fifoOut[40][0];
              muxOutConnector[17] = fifoOut[41][0];
              muxOutConnector[18] = fifoOut[42][0];
              muxOutConnector[19] = fifoOut[43][0];
              muxOutConnector[20] = fifoOut[44][0];
              muxOutConnector[21] = fifoOut[45][0];
              muxOutConnector[22] = fifoOut[46][0];
              muxOutConnector[23] = fifoOut[47][0];
              muxOutConnector[24] = fifoOut[48][0];
              muxOutConnector[25] = fifoOut[49][0];
              muxOutConnector[26] = fifoOut[5][15];
              muxOutConnector[27] = fifoOut[6][15];
              muxOutConnector[28] = fifoOut[7][15];
              muxOutConnector[29] = fifoOut[8][15];
              muxOutConnector[30] = fifoOut[9][15];
              muxOutConnector[31] = fifoOut[10][15];
              muxOutConnector[32] = fifoOut[11][15];
              muxOutConnector[33] = fifoOut[12][15];
              muxOutConnector[34] = fifoOut[13][15];
              muxOutConnector[35] = fifoOut[14][15];
              muxOutConnector[36] = fifoOut[15][15];
              muxOutConnector[37] = fifoOut[16][15];
              muxOutConnector[38] = fifoOut[17][15];
              muxOutConnector[39] = fifoOut[18][15];
              muxOutConnector[40] = fifoOut[19][15];
              muxOutConnector[41] = fifoOut[20][15];
              muxOutConnector[42] = fifoOut[21][15];
              muxOutConnector[43] = fifoOut[22][15];
              muxOutConnector[44] = fifoOut[23][15];
              muxOutConnector[45] = fifoOut[24][15];
              muxOutConnector[46] = fifoOut[25][15];
              muxOutConnector[47] = fifoOut[0][14];
              muxOutConnector[48] = fifoOut[1][14];
              muxOutConnector[49] = fifoOut[2][14];
              muxOutConnector[50] = fifoOut[3][14];
              muxOutConnector[51] = fifoOut[4][14];
         end
         7: begin
              muxOutConnector[0] = fifoOut[50][1];
              muxOutConnector[1] = fifoOut[51][1];
              muxOutConnector[2] = fifoOut[26][0];
              muxOutConnector[3] = fifoOut[27][0];
              muxOutConnector[4] = fifoOut[28][0];
              muxOutConnector[5] = fifoOut[29][0];
              muxOutConnector[6] = fifoOut[30][0];
              muxOutConnector[7] = fifoOut[31][0];
              muxOutConnector[8] = fifoOut[32][0];
              muxOutConnector[9] = fifoOut[33][0];
              muxOutConnector[10] = fifoOut[34][0];
              muxOutConnector[11] = fifoOut[35][0];
              muxOutConnector[12] = fifoOut[36][0];
              muxOutConnector[13] = fifoOut[37][0];
              muxOutConnector[14] = fifoOut[38][0];
              muxOutConnector[15] = fifoOut[39][0];
              muxOutConnector[16] = fifoOut[40][0];
              muxOutConnector[17] = fifoOut[41][0];
              muxOutConnector[18] = fifoOut[42][0];
              muxOutConnector[19] = fifoOut[43][0];
              muxOutConnector[20] = fifoOut[44][0];
              muxOutConnector[21] = fifoOut[45][0];
              muxOutConnector[22] = fifoOut[46][0];
              muxOutConnector[23] = fifoOut[47][0];
              muxOutConnector[24] = fifoOut[48][0];
              muxOutConnector[25] = fifoOut[49][0];
              muxOutConnector[26] = fifoOut[5][15];
              muxOutConnector[27] = fifoOut[6][15];
              muxOutConnector[28] = fifoOut[7][15];
              muxOutConnector[29] = fifoOut[8][15];
              muxOutConnector[30] = fifoOut[9][15];
              muxOutConnector[31] = fifoOut[10][15];
              muxOutConnector[32] = fifoOut[11][15];
              muxOutConnector[33] = fifoOut[12][15];
              muxOutConnector[34] = fifoOut[13][15];
              muxOutConnector[35] = fifoOut[14][15];
              muxOutConnector[36] = fifoOut[15][15];
              muxOutConnector[37] = fifoOut[16][15];
              muxOutConnector[38] = fifoOut[17][15];
              muxOutConnector[39] = fifoOut[18][15];
              muxOutConnector[40] = fifoOut[19][15];
              muxOutConnector[41] = fifoOut[20][15];
              muxOutConnector[42] = fifoOut[21][15];
              muxOutConnector[43] = fifoOut[22][15];
              muxOutConnector[44] = fifoOut[23][15];
              muxOutConnector[45] = fifoOut[24][15];
              muxOutConnector[46] = fifoOut[25][15];
              muxOutConnector[47] = fifoOut[0][14];
              muxOutConnector[48] = fifoOut[1][14];
              muxOutConnector[49] = fifoOut[2][14];
              muxOutConnector[50] = fifoOut[3][14];
              muxOutConnector[51] = fifoOut[4][14];
         end
         8: begin
              muxOutConnector[0] = fifoOut[50][1];
              muxOutConnector[1] = fifoOut[51][1];
              muxOutConnector[2] = fifoOut[26][0];
              muxOutConnector[3] = fifoOut[27][0];
              muxOutConnector[4] = fifoOut[28][0];
              muxOutConnector[5] = fifoOut[29][0];
              muxOutConnector[6] = fifoOut[30][0];
              muxOutConnector[7] = fifoOut[31][0];
              muxOutConnector[8] = fifoOut[32][0];
              muxOutConnector[9] = fifoOut[33][0];
              muxOutConnector[10] = fifoOut[34][0];
              muxOutConnector[11] = fifoOut[35][0];
              muxOutConnector[12] = fifoOut[36][0];
              muxOutConnector[13] = fifoOut[37][0];
              muxOutConnector[14] = fifoOut[38][0];
              muxOutConnector[15] = fifoOut[39][0];
              muxOutConnector[16] = fifoOut[40][0];
              muxOutConnector[17] = fifoOut[41][0];
              muxOutConnector[18] = fifoOut[42][0];
              muxOutConnector[19] = fifoOut[43][0];
              muxOutConnector[20] = fifoOut[44][0];
              muxOutConnector[21] = fifoOut[45][0];
              muxOutConnector[22] = fifoOut[46][0];
              muxOutConnector[23] = fifoOut[47][0];
              muxOutConnector[24] = fifoOut[48][0];
              muxOutConnector[25] = fifoOut[49][0];
              muxOutConnector[26] = fifoOut[5][15];
              muxOutConnector[27] = fifoOut[6][15];
              muxOutConnector[28] = fifoOut[7][15];
              muxOutConnector[29] = fifoOut[8][15];
              muxOutConnector[30] = fifoOut[9][15];
              muxOutConnector[31] = fifoOut[10][15];
              muxOutConnector[32] = fifoOut[11][15];
              muxOutConnector[33] = fifoOut[12][15];
              muxOutConnector[34] = fifoOut[13][15];
              muxOutConnector[35] = fifoOut[14][15];
              muxOutConnector[36] = fifoOut[15][15];
              muxOutConnector[37] = fifoOut[16][15];
              muxOutConnector[38] = fifoOut[17][15];
              muxOutConnector[39] = fifoOut[18][15];
              muxOutConnector[40] = fifoOut[19][15];
              muxOutConnector[41] = fifoOut[20][15];
              muxOutConnector[42] = fifoOut[21][15];
              muxOutConnector[43] = fifoOut[22][15];
              muxOutConnector[44] = fifoOut[23][15];
              muxOutConnector[45] = fifoOut[24][15];
              muxOutConnector[46] = fifoOut[25][15];
              muxOutConnector[47] = fifoOut[0][14];
              muxOutConnector[48] = fifoOut[1][14];
              muxOutConnector[49] = fifoOut[2][14];
              muxOutConnector[50] = fifoOut[3][14];
              muxOutConnector[51] = fifoOut[4][14];
         end
         9: begin
              muxOutConnector[0] = fifoOut[50][1];
              muxOutConnector[1] = fifoOut[51][1];
              muxOutConnector[2] = fifoOut[26][0];
              muxOutConnector[3] = fifoOut[27][0];
              muxOutConnector[4] = fifoOut[28][0];
              muxOutConnector[5] = fifoOut[29][0];
              muxOutConnector[6] = fifoOut[30][0];
              muxOutConnector[7] = fifoOut[31][0];
              muxOutConnector[8] = fifoOut[32][0];
              muxOutConnector[9] = fifoOut[33][0];
              muxOutConnector[10] = fifoOut[34][0];
              muxOutConnector[11] = fifoOut[35][0];
              muxOutConnector[12] = fifoOut[36][0];
              muxOutConnector[13] = fifoOut[37][0];
              muxOutConnector[14] = fifoOut[38][0];
              muxOutConnector[15] = fifoOut[39][0];
              muxOutConnector[16] = fifoOut[40][0];
              muxOutConnector[17] = fifoOut[41][0];
              muxOutConnector[18] = fifoOut[42][0];
              muxOutConnector[19] = fifoOut[43][0];
              muxOutConnector[20] = fifoOut[44][0];
              muxOutConnector[21] = fifoOut[45][0];
              muxOutConnector[22] = fifoOut[46][0];
              muxOutConnector[23] = fifoOut[47][0];
              muxOutConnector[24] = fifoOut[48][0];
              muxOutConnector[25] = fifoOut[49][0];
              muxOutConnector[26] = fifoOut[5][15];
              muxOutConnector[27] = fifoOut[6][15];
              muxOutConnector[28] = fifoOut[7][15];
              muxOutConnector[29] = fifoOut[8][15];
              muxOutConnector[30] = fifoOut[9][15];
              muxOutConnector[31] = fifoOut[10][15];
              muxOutConnector[32] = fifoOut[11][15];
              muxOutConnector[33] = fifoOut[12][15];
              muxOutConnector[34] = fifoOut[13][15];
              muxOutConnector[35] = fifoOut[14][15];
              muxOutConnector[36] = fifoOut[15][15];
              muxOutConnector[37] = fifoOut[16][15];
              muxOutConnector[38] = fifoOut[17][15];
              muxOutConnector[39] = fifoOut[18][15];
              muxOutConnector[40] = fifoOut[19][15];
              muxOutConnector[41] = fifoOut[20][15];
              muxOutConnector[42] = fifoOut[21][15];
              muxOutConnector[43] = fifoOut[22][15];
              muxOutConnector[44] = fifoOut[23][15];
              muxOutConnector[45] = fifoOut[24][15];
              muxOutConnector[46] = fifoOut[25][15];
              muxOutConnector[47] = fifoOut[0][14];
              muxOutConnector[48] = fifoOut[1][14];
              muxOutConnector[49] = fifoOut[2][14];
              muxOutConnector[50] = fifoOut[3][14];
              muxOutConnector[51] = fifoOut[4][14];
         end
         10: begin
              muxOutConnector[0] = fifoOut[50][1];
              muxOutConnector[1] = fifoOut[51][1];
              muxOutConnector[2] = fifoOut[26][0];
              muxOutConnector[3] = fifoOut[27][0];
              muxOutConnector[4] = fifoOut[28][0];
              muxOutConnector[5] = fifoOut[29][0];
              muxOutConnector[6] = fifoOut[30][0];
              muxOutConnector[7] = fifoOut[31][0];
              muxOutConnector[8] = fifoOut[32][0];
              muxOutConnector[9] = fifoOut[33][0];
              muxOutConnector[10] = fifoOut[34][0];
              muxOutConnector[11] = fifoOut[35][0];
              muxOutConnector[12] = fifoOut[36][0];
              muxOutConnector[13] = fifoOut[37][0];
              muxOutConnector[14] = fifoOut[0][6];
              muxOutConnector[15] = fifoOut[1][6];
              muxOutConnector[16] = fifoOut[2][6];
              muxOutConnector[17] = fifoOut[3][6];
              muxOutConnector[18] = fifoOut[4][6];
              muxOutConnector[19] = fifoOut[5][6];
              muxOutConnector[20] = fifoOut[6][6];
              muxOutConnector[21] = fifoOut[7][6];
              muxOutConnector[22] = fifoOut[8][6];
              muxOutConnector[23] = fifoOut[9][6];
              muxOutConnector[24] = fifoOut[10][6];
              muxOutConnector[25] = fifoOut[11][6];
              muxOutConnector[26] = fifoOut[5][15];
              muxOutConnector[27] = fifoOut[6][15];
              muxOutConnector[28] = fifoOut[7][15];
              muxOutConnector[29] = fifoOut[8][15];
              muxOutConnector[30] = fifoOut[9][15];
              muxOutConnector[31] = fifoOut[10][15];
              muxOutConnector[32] = fifoOut[11][15];
              muxOutConnector[33] = fifoOut[12][15];
              muxOutConnector[34] = fifoOut[13][15];
              muxOutConnector[35] = fifoOut[14][15];
              muxOutConnector[36] = fifoOut[15][15];
              muxOutConnector[37] = fifoOut[16][15];
              muxOutConnector[38] = fifoOut[17][15];
              muxOutConnector[39] = fifoOut[18][15];
              muxOutConnector[40] = fifoOut[19][15];
              muxOutConnector[41] = fifoOut[20][15];
              muxOutConnector[42] = fifoOut[21][15];
              muxOutConnector[43] = fifoOut[22][15];
              muxOutConnector[44] = fifoOut[23][15];
              muxOutConnector[45] = fifoOut[24][15];
              muxOutConnector[46] = fifoOut[25][15];
              muxOutConnector[47] = fifoOut[0][14];
              muxOutConnector[48] = fifoOut[1][14];
              muxOutConnector[49] = fifoOut[2][14];
              muxOutConnector[50] = fifoOut[3][14];
              muxOutConnector[51] = fifoOut[4][14];
         end
         11: begin
              muxOutConnector[0] = fifoOut[12][7];
              muxOutConnector[1] = fifoOut[13][7];
              muxOutConnector[2] = fifoOut[14][7];
              muxOutConnector[3] = fifoOut[15][7];
              muxOutConnector[4] = fifoOut[16][7];
              muxOutConnector[5] = fifoOut[17][7];
              muxOutConnector[6] = fifoOut[18][7];
              muxOutConnector[7] = fifoOut[19][7];
              muxOutConnector[8] = fifoOut[20][7];
              muxOutConnector[9] = fifoOut[21][7];
              muxOutConnector[10] = fifoOut[22][7];
              muxOutConnector[11] = fifoOut[23][7];
              muxOutConnector[12] = fifoOut[24][7];
              muxOutConnector[13] = fifoOut[25][7];
              muxOutConnector[14] = fifoOut[0][6];
              muxOutConnector[15] = fifoOut[1][6];
              muxOutConnector[16] = fifoOut[2][6];
              muxOutConnector[17] = fifoOut[3][6];
              muxOutConnector[18] = fifoOut[4][6];
              muxOutConnector[19] = fifoOut[5][6];
              muxOutConnector[20] = fifoOut[6][6];
              muxOutConnector[21] = fifoOut[7][6];
              muxOutConnector[22] = fifoOut[8][6];
              muxOutConnector[23] = fifoOut[9][6];
              muxOutConnector[24] = fifoOut[10][6];
              muxOutConnector[25] = fifoOut[11][6];
              muxOutConnector[26] = fifoOut[5][15];
              muxOutConnector[27] = fifoOut[6][15];
              muxOutConnector[28] = fifoOut[7][15];
              muxOutConnector[29] = fifoOut[8][15];
              muxOutConnector[30] = fifoOut[9][15];
              muxOutConnector[31] = fifoOut[10][15];
              muxOutConnector[32] = fifoOut[11][15];
              muxOutConnector[33] = fifoOut[12][15];
              muxOutConnector[34] = fifoOut[13][15];
              muxOutConnector[35] = fifoOut[14][15];
              muxOutConnector[36] = fifoOut[15][15];
              muxOutConnector[37] = fifoOut[16][15];
              muxOutConnector[38] = fifoOut[17][15];
              muxOutConnector[39] = fifoOut[18][15];
              muxOutConnector[40] = fifoOut[19][15];
              muxOutConnector[41] = fifoOut[20][15];
              muxOutConnector[42] = fifoOut[21][15];
              muxOutConnector[43] = fifoOut[22][15];
              muxOutConnector[44] = fifoOut[23][15];
              muxOutConnector[45] = fifoOut[24][15];
              muxOutConnector[46] = fifoOut[25][15];
              muxOutConnector[47] = fifoOut[0][14];
              muxOutConnector[48] = fifoOut[1][14];
              muxOutConnector[49] = fifoOut[2][14];
              muxOutConnector[50] = fifoOut[3][14];
              muxOutConnector[51] = fifoOut[4][14];
         end
         12: begin
              muxOutConnector[0] = fifoOut[12][7];
              muxOutConnector[1] = fifoOut[13][7];
              muxOutConnector[2] = fifoOut[14][7];
              muxOutConnector[3] = fifoOut[15][7];
              muxOutConnector[4] = fifoOut[16][7];
              muxOutConnector[5] = fifoOut[17][7];
              muxOutConnector[6] = fifoOut[18][7];
              muxOutConnector[7] = fifoOut[19][7];
              muxOutConnector[8] = fifoOut[20][7];
              muxOutConnector[9] = fifoOut[21][7];
              muxOutConnector[10] = fifoOut[22][7];
              muxOutConnector[11] = fifoOut[23][7];
              muxOutConnector[12] = fifoOut[24][7];
              muxOutConnector[13] = fifoOut[25][7];
              muxOutConnector[14] = fifoOut[0][6];
              muxOutConnector[15] = fifoOut[1][6];
              muxOutConnector[16] = fifoOut[2][6];
              muxOutConnector[17] = fifoOut[3][6];
              muxOutConnector[18] = fifoOut[4][6];
              muxOutConnector[19] = fifoOut[5][6];
              muxOutConnector[20] = fifoOut[6][6];
              muxOutConnector[21] = fifoOut[7][6];
              muxOutConnector[22] = fifoOut[8][6];
              muxOutConnector[23] = fifoOut[9][6];
              muxOutConnector[24] = fifoOut[10][6];
              muxOutConnector[25] = fifoOut[11][6];
              muxOutConnector[26] = fifoOut[5][15];
              muxOutConnector[27] = fifoOut[6][15];
              muxOutConnector[28] = fifoOut[7][15];
              muxOutConnector[29] = fifoOut[8][15];
              muxOutConnector[30] = fifoOut[9][15];
              muxOutConnector[31] = fifoOut[10][15];
              muxOutConnector[32] = fifoOut[11][15];
              muxOutConnector[33] = fifoOut[12][15];
              muxOutConnector[34] = fifoOut[13][15];
              muxOutConnector[35] = fifoOut[14][15];
              muxOutConnector[36] = fifoOut[15][15];
              muxOutConnector[37] = fifoOut[16][15];
              muxOutConnector[38] = fifoOut[17][15];
              muxOutConnector[39] = fifoOut[18][15];
              muxOutConnector[40] = fifoOut[19][15];
              muxOutConnector[41] = fifoOut[20][15];
              muxOutConnector[42] = fifoOut[21][15];
              muxOutConnector[43] = fifoOut[22][15];
              muxOutConnector[44] = fifoOut[23][15];
              muxOutConnector[45] = fifoOut[24][15];
              muxOutConnector[46] = fifoOut[25][15];
              muxOutConnector[47] = fifoOut[0][14];
              muxOutConnector[48] = fifoOut[1][14];
              muxOutConnector[49] = fifoOut[2][14];
              muxOutConnector[50] = fifoOut[3][14];
              muxOutConnector[51] = fifoOut[4][14];
         end
         13: begin
              muxOutConnector[0] = fifoOut[12][7];
              muxOutConnector[1] = fifoOut[13][7];
              muxOutConnector[2] = fifoOut[14][7];
              muxOutConnector[3] = fifoOut[15][7];
              muxOutConnector[4] = fifoOut[16][7];
              muxOutConnector[5] = fifoOut[17][7];
              muxOutConnector[6] = fifoOut[18][7];
              muxOutConnector[7] = fifoOut[19][7];
              muxOutConnector[8] = fifoOut[20][7];
              muxOutConnector[9] = fifoOut[21][7];
              muxOutConnector[10] = fifoOut[22][7];
              muxOutConnector[11] = fifoOut[23][7];
              muxOutConnector[12] = fifoOut[24][7];
              muxOutConnector[13] = fifoOut[25][7];
              muxOutConnector[14] = fifoOut[0][6];
              muxOutConnector[15] = fifoOut[1][6];
              muxOutConnector[16] = fifoOut[2][6];
              muxOutConnector[17] = fifoOut[3][6];
              muxOutConnector[18] = fifoOut[4][6];
              muxOutConnector[19] = fifoOut[5][6];
              muxOutConnector[20] = fifoOut[6][6];
              muxOutConnector[21] = fifoOut[7][6];
              muxOutConnector[22] = fifoOut[8][6];
              muxOutConnector[23] = fifoOut[9][6];
              muxOutConnector[24] = fifoOut[10][6];
              muxOutConnector[25] = fifoOut[11][6];
              muxOutConnector[26] = fifoOut[5][15];
              muxOutConnector[27] = fifoOut[6][15];
              muxOutConnector[28] = fifoOut[7][15];
              muxOutConnector[29] = fifoOut[8][15];
              muxOutConnector[30] = fifoOut[9][15];
              muxOutConnector[31] = fifoOut[10][15];
              muxOutConnector[32] = fifoOut[11][15];
              muxOutConnector[33] = fifoOut[12][15];
              muxOutConnector[34] = fifoOut[13][15];
              muxOutConnector[35] = fifoOut[14][15];
              muxOutConnector[36] = fifoOut[15][15];
              muxOutConnector[37] = fifoOut[16][15];
              muxOutConnector[38] = fifoOut[17][15];
              muxOutConnector[39] = fifoOut[18][15];
              muxOutConnector[40] = fifoOut[19][15];
              muxOutConnector[41] = fifoOut[20][15];
              muxOutConnector[42] = fifoOut[21][15];
              muxOutConnector[43] = fifoOut[22][15];
              muxOutConnector[44] = fifoOut[23][15];
              muxOutConnector[45] = fifoOut[24][15];
              muxOutConnector[46] = fifoOut[25][15];
              muxOutConnector[47] = fifoOut[0][14];
              muxOutConnector[48] = fifoOut[1][14];
              muxOutConnector[49] = fifoOut[2][14];
              muxOutConnector[50] = fifoOut[3][14];
              muxOutConnector[51] = fifoOut[4][14];
         end
         14: begin
              muxOutConnector[0] = fifoOut[12][7];
              muxOutConnector[1] = fifoOut[13][7];
              muxOutConnector[2] = fifoOut[14][7];
              muxOutConnector[3] = fifoOut[15][7];
              muxOutConnector[4] = fifoOut[16][7];
              muxOutConnector[5] = fifoOut[17][7];
              muxOutConnector[6] = fifoOut[18][7];
              muxOutConnector[7] = fifoOut[19][7];
              muxOutConnector[8] = fifoOut[20][7];
              muxOutConnector[9] = fifoOut[21][7];
              muxOutConnector[10] = fifoOut[22][7];
              muxOutConnector[11] = fifoOut[23][7];
              muxOutConnector[12] = fifoOut[24][7];
              muxOutConnector[13] = fifoOut[25][7];
              muxOutConnector[14] = fifoOut[0][6];
              muxOutConnector[15] = fifoOut[1][6];
              muxOutConnector[16] = fifoOut[2][6];
              muxOutConnector[17] = fifoOut[3][6];
              muxOutConnector[18] = fifoOut[4][6];
              muxOutConnector[19] = fifoOut[5][6];
              muxOutConnector[20] = fifoOut[6][6];
              muxOutConnector[21] = fifoOut[7][6];
              muxOutConnector[22] = fifoOut[8][6];
              muxOutConnector[23] = fifoOut[9][6];
              muxOutConnector[24] = fifoOut[10][6];
              muxOutConnector[25] = fifoOut[11][6];
              muxOutConnector[26] = fifoOut[5][15];
              muxOutConnector[27] = fifoOut[6][15];
              muxOutConnector[28] = fifoOut[7][15];
              muxOutConnector[29] = fifoOut[8][15];
              muxOutConnector[30] = fifoOut[9][15];
              muxOutConnector[31] = fifoOut[10][15];
              muxOutConnector[32] = fifoOut[11][15];
              muxOutConnector[33] = fifoOut[12][15];
              muxOutConnector[34] = fifoOut[13][15];
              muxOutConnector[35] = fifoOut[14][15];
              muxOutConnector[36] = fifoOut[15][15];
              muxOutConnector[37] = fifoOut[16][15];
              muxOutConnector[38] = fifoOut[17][15];
              muxOutConnector[39] = fifoOut[18][15];
              muxOutConnector[40] = fifoOut[19][15];
              muxOutConnector[41] = fifoOut[20][15];
              muxOutConnector[42] = fifoOut[21][15];
              muxOutConnector[43] = fifoOut[22][15];
              muxOutConnector[44] = fifoOut[23][15];
              muxOutConnector[45] = fifoOut[24][15];
              muxOutConnector[46] = fifoOut[25][15];
              muxOutConnector[47] = fifoOut[0][14];
              muxOutConnector[48] = fifoOut[1][14];
              muxOutConnector[49] = fifoOut[2][14];
              muxOutConnector[50] = fifoOut[3][14];
              muxOutConnector[51] = fifoOut[4][14];
         end
         15: begin
              muxOutConnector[0] = fifoOut[12][7];
              muxOutConnector[1] = fifoOut[13][7];
              muxOutConnector[2] = fifoOut[14][7];
              muxOutConnector[3] = fifoOut[15][7];
              muxOutConnector[4] = fifoOut[16][7];
              muxOutConnector[5] = fifoOut[17][7];
              muxOutConnector[6] = fifoOut[18][7];
              muxOutConnector[7] = fifoOut[19][7];
              muxOutConnector[8] = fifoOut[20][7];
              muxOutConnector[9] = fifoOut[21][7];
              muxOutConnector[10] = fifoOut[22][7];
              muxOutConnector[11] = fifoOut[23][7];
              muxOutConnector[12] = fifoOut[24][7];
              muxOutConnector[13] = fifoOut[25][7];
              muxOutConnector[14] = fifoOut[0][6];
              muxOutConnector[15] = fifoOut[1][6];
              muxOutConnector[16] = fifoOut[2][6];
              muxOutConnector[17] = fifoOut[3][6];
              muxOutConnector[18] = fifoOut[4][6];
              muxOutConnector[19] = fifoOut[5][6];
              muxOutConnector[20] = fifoOut[6][6];
              muxOutConnector[21] = fifoOut[7][6];
              muxOutConnector[22] = fifoOut[8][6];
              muxOutConnector[23] = fifoOut[9][6];
              muxOutConnector[24] = fifoOut[10][6];
              muxOutConnector[25] = fifoOut[11][6];
              muxOutConnector[26] = fifoOut[5][15];
              muxOutConnector[27] = fifoOut[6][15];
              muxOutConnector[28] = fifoOut[7][15];
              muxOutConnector[29] = fifoOut[8][15];
              muxOutConnector[30] = fifoOut[9][15];
              muxOutConnector[31] = fifoOut[10][15];
              muxOutConnector[32] = fifoOut[11][15];
              muxOutConnector[33] = fifoOut[12][15];
              muxOutConnector[34] = fifoOut[13][15];
              muxOutConnector[35] = fifoOut[14][15];
              muxOutConnector[36] = fifoOut[15][15];
              muxOutConnector[37] = fifoOut[16][15];
              muxOutConnector[38] = fifoOut[38][11];
              muxOutConnector[39] = fifoOut[39][11];
              muxOutConnector[40] = fifoOut[40][11];
              muxOutConnector[41] = fifoOut[41][11];
              muxOutConnector[42] = fifoOut[42][11];
              muxOutConnector[43] = fifoOut[43][11];
              muxOutConnector[44] = fifoOut[44][11];
              muxOutConnector[45] = fifoOut[45][11];
              muxOutConnector[46] = fifoOut[46][11];
              muxOutConnector[47] = fifoOut[47][11];
              muxOutConnector[48] = fifoOut[48][11];
              muxOutConnector[49] = fifoOut[49][11];
              muxOutConnector[50] = fifoOut[50][11];
              muxOutConnector[51] = fifoOut[51][11];
         end
         16: begin
              muxOutConnector[0] = fifoOut[12][7];
              muxOutConnector[1] = fifoOut[13][7];
              muxOutConnector[2] = fifoOut[14][7];
              muxOutConnector[3] = fifoOut[15][7];
              muxOutConnector[4] = fifoOut[16][7];
              muxOutConnector[5] = fifoOut[17][7];
              muxOutConnector[6] = fifoOut[18][7];
              muxOutConnector[7] = fifoOut[19][7];
              muxOutConnector[8] = fifoOut[20][7];
              muxOutConnector[9] = fifoOut[21][7];
              muxOutConnector[10] = fifoOut[22][7];
              muxOutConnector[11] = fifoOut[23][7];
              muxOutConnector[12] = fifoOut[24][7];
              muxOutConnector[13] = fifoOut[25][7];
              muxOutConnector[14] = fifoOut[0][6];
              muxOutConnector[15] = fifoOut[1][6];
              muxOutConnector[16] = fifoOut[2][6];
              muxOutConnector[17] = fifoOut[3][6];
              muxOutConnector[18] = fifoOut[4][6];
              muxOutConnector[19] = fifoOut[5][6];
              muxOutConnector[20] = fifoOut[6][6];
              muxOutConnector[21] = fifoOut[7][6];
              muxOutConnector[22] = fifoOut[8][6];
              muxOutConnector[23] = fifoOut[9][6];
              muxOutConnector[24] = fifoOut[10][6];
              muxOutConnector[25] = fifoOut[11][6];
              muxOutConnector[26] = fifoOut[26][11];
              muxOutConnector[27] = fifoOut[27][11];
              muxOutConnector[28] = fifoOut[28][11];
              muxOutConnector[29] = fifoOut[29][11];
              muxOutConnector[30] = fifoOut[30][11];
              muxOutConnector[31] = fifoOut[31][11];
              muxOutConnector[32] = fifoOut[32][11];
              muxOutConnector[33] = fifoOut[33][11];
              muxOutConnector[34] = fifoOut[34][11];
              muxOutConnector[35] = fifoOut[35][11];
              muxOutConnector[36] = fifoOut[36][11];
              muxOutConnector[37] = fifoOut[37][11];
              muxOutConnector[38] = fifoOut[38][11];
              muxOutConnector[39] = fifoOut[39][11];
              muxOutConnector[40] = fifoOut[40][11];
              muxOutConnector[41] = fifoOut[41][11];
              muxOutConnector[42] = fifoOut[42][11];
              muxOutConnector[43] = fifoOut[43][11];
              muxOutConnector[44] = fifoOut[44][11];
              muxOutConnector[45] = fifoOut[45][11];
              muxOutConnector[46] = fifoOut[46][11];
              muxOutConnector[47] = fifoOut[47][11];
              muxOutConnector[48] = fifoOut[48][11];
              muxOutConnector[49] = fifoOut[49][11];
              muxOutConnector[50] = fifoOut[50][11];
              muxOutConnector[51] = fifoOut[51][11];
         end
         17: begin
              muxOutConnector[0] = fifoOut[12][7];
              muxOutConnector[1] = fifoOut[13][7];
              muxOutConnector[2] = fifoOut[14][7];
              muxOutConnector[3] = fifoOut[15][7];
              muxOutConnector[4] = fifoOut[16][7];
              muxOutConnector[5] = fifoOut[17][7];
              muxOutConnector[6] = fifoOut[18][7];
              muxOutConnector[7] = fifoOut[19][7];
              muxOutConnector[8] = fifoOut[20][7];
              muxOutConnector[9] = fifoOut[21][7];
              muxOutConnector[10] = fifoOut[22][7];
              muxOutConnector[11] = fifoOut[23][7];
              muxOutConnector[12] = fifoOut[24][7];
              muxOutConnector[13] = fifoOut[25][7];
              muxOutConnector[14] = fifoOut[0][6];
              muxOutConnector[15] = fifoOut[1][6];
              muxOutConnector[16] = fifoOut[2][6];
              muxOutConnector[17] = fifoOut[3][6];
              muxOutConnector[18] = fifoOut[4][6];
              muxOutConnector[19] = fifoOut[5][6];
              muxOutConnector[20] = fifoOut[6][6];
              muxOutConnector[21] = fifoOut[7][6];
              muxOutConnector[22] = fifoOut[8][6];
              muxOutConnector[23] = fifoOut[9][6];
              muxOutConnector[24] = fifoOut[10][6];
              muxOutConnector[25] = fifoOut[11][6];
              muxOutConnector[26] = fifoOut[26][11];
              muxOutConnector[27] = fifoOut[27][11];
              muxOutConnector[28] = fifoOut[28][11];
              muxOutConnector[29] = fifoOut[29][11];
              muxOutConnector[30] = fifoOut[30][11];
              muxOutConnector[31] = fifoOut[31][11];
              muxOutConnector[32] = fifoOut[32][11];
              muxOutConnector[33] = fifoOut[33][11];
              muxOutConnector[34] = fifoOut[34][11];
              muxOutConnector[35] = fifoOut[35][11];
              muxOutConnector[36] = fifoOut[36][11];
              muxOutConnector[37] = fifoOut[37][11];
              muxOutConnector[38] = fifoOut[38][11];
              muxOutConnector[39] = fifoOut[39][11];
              muxOutConnector[40] = fifoOut[40][11];
              muxOutConnector[41] = fifoOut[41][11];
              muxOutConnector[42] = fifoOut[42][11];
              muxOutConnector[43] = fifoOut[43][11];
              muxOutConnector[44] = fifoOut[44][11];
              muxOutConnector[45] = fifoOut[45][11];
              muxOutConnector[46] = fifoOut[46][11];
              muxOutConnector[47] = fifoOut[47][11];
              muxOutConnector[48] = fifoOut[48][11];
              muxOutConnector[49] = fifoOut[49][11];
              muxOutConnector[50] = fifoOut[50][11];
              muxOutConnector[51] = fifoOut[51][11];
         end
         18: begin
              muxOutConnector[0] = fifoOut[12][7];
              muxOutConnector[1] = fifoOut[13][7];
              muxOutConnector[2] = fifoOut[14][7];
              muxOutConnector[3] = fifoOut[15][7];
              muxOutConnector[4] = fifoOut[16][7];
              muxOutConnector[5] = fifoOut[17][7];
              muxOutConnector[6] = fifoOut[18][7];
              muxOutConnector[7] = fifoOut[19][7];
              muxOutConnector[8] = fifoOut[20][7];
              muxOutConnector[9] = fifoOut[21][7];
              muxOutConnector[10] = fifoOut[22][7];
              muxOutConnector[11] = fifoOut[23][7];
              muxOutConnector[12] = fifoOut[24][7];
              muxOutConnector[13] = fifoOut[25][7];
              muxOutConnector[14] = fifoOut[0][6];
              muxOutConnector[15] = fifoOut[1][6];
              muxOutConnector[16] = fifoOut[2][6];
              muxOutConnector[17] = fifoOut[3][6];
              muxOutConnector[18] = fifoOut[4][6];
              muxOutConnector[19] = fifoOut[5][6];
              muxOutConnector[20] = fifoOut[6][6];
              muxOutConnector[21] = fifoOut[7][6];
              muxOutConnector[22] = fifoOut[8][6];
              muxOutConnector[23] = fifoOut[9][6];
              muxOutConnector[24] = fifoOut[10][6];
              muxOutConnector[25] = fifoOut[11][6];
              muxOutConnector[26] = fifoOut[26][11];
              muxOutConnector[27] = fifoOut[27][11];
              muxOutConnector[28] = fifoOut[28][11];
              muxOutConnector[29] = fifoOut[29][11];
              muxOutConnector[30] = fifoOut[30][11];
              muxOutConnector[31] = fifoOut[31][11];
              muxOutConnector[32] = fifoOut[32][11];
              muxOutConnector[33] = fifoOut[33][11];
              muxOutConnector[34] = fifoOut[34][11];
              muxOutConnector[35] = fifoOut[35][11];
              muxOutConnector[36] = fifoOut[36][11];
              muxOutConnector[37] = fifoOut[37][11];
              muxOutConnector[38] = fifoOut[38][11];
              muxOutConnector[39] = fifoOut[39][11];
              muxOutConnector[40] = fifoOut[40][11];
              muxOutConnector[41] = fifoOut[41][11];
              muxOutConnector[42] = fifoOut[42][11];
              muxOutConnector[43] = fifoOut[43][11];
              muxOutConnector[44] = fifoOut[44][11];
              muxOutConnector[45] = fifoOut[45][11];
              muxOutConnector[46] = fifoOut[46][11];
              muxOutConnector[47] = fifoOut[47][11];
              muxOutConnector[48] = fifoOut[48][11];
              muxOutConnector[49] = fifoOut[49][11];
              muxOutConnector[50] = fifoOut[50][11];
              muxOutConnector[51] = fifoOut[51][11];
         end
         19: begin
              muxOutConnector[0] = fifoOut[12][7];
              muxOutConnector[1] = fifoOut[13][7];
              muxOutConnector[2] = fifoOut[14][7];
              muxOutConnector[3] = fifoOut[15][7];
              muxOutConnector[4] = fifoOut[16][7];
              muxOutConnector[5] = fifoOut[17][7];
              muxOutConnector[6] = fifoOut[18][7];
              muxOutConnector[7] = fifoOut[19][7];
              muxOutConnector[8] = fifoOut[20][7];
              muxOutConnector[9] = fifoOut[21][7];
              muxOutConnector[10] = fifoOut[22][7];
              muxOutConnector[11] = fifoOut[23][7];
              muxOutConnector[12] = fifoOut[24][7];
              muxOutConnector[13] = fifoOut[25][7];
              muxOutConnector[14] = fifoOut[0][6];
              muxOutConnector[15] = fifoOut[1][6];
              muxOutConnector[16] = fifoOut[2][6];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[26][11];
              muxOutConnector[27] = fifoOut[27][11];
              muxOutConnector[28] = fifoOut[28][11];
              muxOutConnector[29] = fifoOut[29][11];
              muxOutConnector[30] = fifoOut[30][11];
              muxOutConnector[31] = fifoOut[31][11];
              muxOutConnector[32] = fifoOut[32][11];
              muxOutConnector[33] = fifoOut[33][11];
              muxOutConnector[34] = fifoOut[34][11];
              muxOutConnector[35] = fifoOut[35][11];
              muxOutConnector[36] = fifoOut[36][11];
              muxOutConnector[37] = fifoOut[37][11];
              muxOutConnector[38] = fifoOut[38][11];
              muxOutConnector[39] = fifoOut[39][11];
              muxOutConnector[40] = fifoOut[40][11];
              muxOutConnector[41] = fifoOut[41][11];
              muxOutConnector[42] = fifoOut[42][11];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
         end
         default: begin
               for(i=0;i<muxOutSymbols;i=i+1)begin
                muxOutConnector[i] = 0;
              end
         end
//hgjhgbuiguigbigbgbgbui
         endcase
    end
endcase
             end
        endmodule