`timescale 1ns / 1ps
module LMem0To1_511_circ1_ys_scripted(
        muxOut,
        ly0In,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 12;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

reg   feedback_en;
reg [ w - 1 : 0 ]column_1[ r - 1 : 0 ];
reg chip_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(chip_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= column_1[i];
         end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
  feedback_en=rd_en;
      if(wr_en)begin
        chip_en=wr_en;
      end
      else begin
        chip_en=feedback_en;
      end
   if(feedback_en)begin
      for(i = r-1; i > -1; i=i-1) begin
        column_1[i] = fifoOut[i][c-1];
      end
   end
   else begin
      for(i = r-1; i > -1; i=i-1) begin
        column_1[i] = ly0InConnector[i];
      end
    end
end
always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[38][4];
              muxOutConnector[1] = fifoOut[39][4];
              muxOutConnector[2] = fifoOut[40][4];
              muxOutConnector[3] = fifoOut[41][4];
              muxOutConnector[4] = fifoOut[42][4];
              muxOutConnector[5] = fifoOut[43][4];
              muxOutConnector[6] = fifoOut[44][4];
              muxOutConnector[7] = fifoOut[45][4];
              muxOutConnector[8] = fifoOut[46][4];
              muxOutConnector[9] = fifoOut[47][4];
              muxOutConnector[10] = fifoOut[48][4];
              muxOutConnector[11] = fifoOut[49][4];
              muxOutConnector[12] = fifoOut[50][4];
              muxOutConnector[13] = fifoOut[51][4];
              muxOutConnector[14] = fifoOut[26][3];
              muxOutConnector[15] = fifoOut[27][3];
              muxOutConnector[16] = fifoOut[28][3];
              muxOutConnector[17] = fifoOut[29][3];
              muxOutConnector[18] = fifoOut[30][3];
              muxOutConnector[19] = fifoOut[31][3];
              muxOutConnector[20] = fifoOut[32][3];
              muxOutConnector[21] = fifoOut[33][3];
              muxOutConnector[22] = fifoOut[34][3];
              muxOutConnector[23] = fifoOut[35][3];
              muxOutConnector[24] = fifoOut[36][3];
              muxOutConnector[25] = fifoOut[37][3];
              muxOutConnector[26] = fifoOut[26][10];
              muxOutConnector[27] = fifoOut[27][10];
              muxOutConnector[28] = fifoOut[28][10];
              muxOutConnector[29] = fifoOut[29][10];
              muxOutConnector[30] = fifoOut[30][10];
              muxOutConnector[31] = fifoOut[31][10];
              muxOutConnector[32] = fifoOut[32][10];
              muxOutConnector[33] = fifoOut[33][10];
              muxOutConnector[34] = fifoOut[34][10];
              muxOutConnector[35] = fifoOut[35][10];
              muxOutConnector[36] = fifoOut[36][10];
              muxOutConnector[37] = fifoOut[37][10];
              muxOutConnector[38] = fifoOut[38][10];
              muxOutConnector[39] = fifoOut[39][10];
              muxOutConnector[40] = fifoOut[40][10];
              muxOutConnector[41] = fifoOut[41][10];
              muxOutConnector[42] = fifoOut[42][10];
              muxOutConnector[43] = fifoOut[43][10];
              muxOutConnector[44] = fifoOut[44][10];
              muxOutConnector[45] = fifoOut[45][10];
              muxOutConnector[46] = fifoOut[46][10];
              muxOutConnector[47] = fifoOut[47][10];
              muxOutConnector[48] = fifoOut[48][10];
              muxOutConnector[49] = fifoOut[49][10];
              muxOutConnector[50] = fifoOut[50][10];
              muxOutConnector[51] = fifoOut[51][10];
       end
       1: begin
              muxOutConnector[0] = fifoOut[38][4];
              muxOutConnector[1] = fifoOut[39][4];
              muxOutConnector[2] = fifoOut[40][4];
              muxOutConnector[3] = fifoOut[41][4];
              muxOutConnector[4] = fifoOut[42][4];
              muxOutConnector[5] = fifoOut[43][4];
              muxOutConnector[6] = fifoOut[44][4];
              muxOutConnector[7] = fifoOut[45][4];
              muxOutConnector[8] = fifoOut[46][4];
              muxOutConnector[9] = fifoOut[47][4];
              muxOutConnector[10] = fifoOut[48][4];
              muxOutConnector[11] = fifoOut[49][4];
              muxOutConnector[12] = fifoOut[50][4];
              muxOutConnector[13] = fifoOut[51][4];
              muxOutConnector[14] = fifoOut[26][3];
              muxOutConnector[15] = fifoOut[27][3];
              muxOutConnector[16] = fifoOut[28][3];
              muxOutConnector[17] = fifoOut[29][3];
              muxOutConnector[18] = fifoOut[30][3];
              muxOutConnector[19] = fifoOut[31][3];
              muxOutConnector[20] = fifoOut[32][3];
              muxOutConnector[21] = fifoOut[33][3];
              muxOutConnector[22] = fifoOut[34][3];
              muxOutConnector[23] = fifoOut[35][3];
              muxOutConnector[24] = fifoOut[36][3];
              muxOutConnector[25] = fifoOut[37][3];
              muxOutConnector[26] = fifoOut[26][10];
              muxOutConnector[27] = fifoOut[27][10];
              muxOutConnector[28] = fifoOut[28][10];
              muxOutConnector[29] = fifoOut[29][10];
              muxOutConnector[30] = fifoOut[30][10];
              muxOutConnector[31] = fifoOut[31][10];
              muxOutConnector[32] = fifoOut[32][10];
              muxOutConnector[33] = fifoOut[33][10];
              muxOutConnector[34] = fifoOut[34][10];
              muxOutConnector[35] = fifoOut[35][10];
              muxOutConnector[36] = fifoOut[36][10];
              muxOutConnector[37] = fifoOut[37][10];
              muxOutConnector[38] = fifoOut[38][10];
              muxOutConnector[39] = fifoOut[39][10];
              muxOutConnector[40] = fifoOut[40][10];
              muxOutConnector[41] = fifoOut[41][10];
              muxOutConnector[42] = fifoOut[42][10];
              muxOutConnector[43] = fifoOut[43][10];
              muxOutConnector[44] = fifoOut[44][10];
              muxOutConnector[45] = fifoOut[45][10];
              muxOutConnector[46] = fifoOut[46][10];
              muxOutConnector[47] = fifoOut[47][10];
              muxOutConnector[48] = fifoOut[48][10];
              muxOutConnector[49] = fifoOut[49][10];
              muxOutConnector[50] = fifoOut[50][10];
              muxOutConnector[51] = fifoOut[51][10];
       end
       2: begin
              muxOutConnector[0] = fifoOut[38][4];
              muxOutConnector[1] = fifoOut[39][4];
              muxOutConnector[2] = fifoOut[40][4];
              muxOutConnector[3] = fifoOut[41][4];
              muxOutConnector[4] = fifoOut[42][4];
              muxOutConnector[5] = fifoOut[43][4];
              muxOutConnector[6] = fifoOut[44][4];
              muxOutConnector[7] = fifoOut[45][4];
              muxOutConnector[8] = fifoOut[46][4];
              muxOutConnector[9] = fifoOut[47][4];
              muxOutConnector[10] = fifoOut[48][4];
              muxOutConnector[11] = fifoOut[49][4];
              muxOutConnector[12] = fifoOut[50][4];
              muxOutConnector[13] = fifoOut[51][4];
              muxOutConnector[14] = fifoOut[26][3];
              muxOutConnector[15] = fifoOut[27][3];
              muxOutConnector[16] = fifoOut[28][3];
              muxOutConnector[17] = fifoOut[29][3];
              muxOutConnector[18] = fifoOut[30][3];
              muxOutConnector[19] = fifoOut[31][3];
              muxOutConnector[20] = fifoOut[32][3];
              muxOutConnector[21] = fifoOut[33][3];
              muxOutConnector[22] = fifoOut[34][3];
              muxOutConnector[23] = fifoOut[35][3];
              muxOutConnector[24] = fifoOut[36][3];
              muxOutConnector[25] = fifoOut[37][3];
              muxOutConnector[26] = fifoOut[26][10];
              muxOutConnector[27] = fifoOut[27][10];
              muxOutConnector[28] = fifoOut[28][10];
              muxOutConnector[29] = fifoOut[29][10];
              muxOutConnector[30] = fifoOut[30][10];
              muxOutConnector[31] = fifoOut[31][10];
              muxOutConnector[32] = fifoOut[32][10];
              muxOutConnector[33] = fifoOut[33][10];
              muxOutConnector[34] = fifoOut[34][10];
              muxOutConnector[35] = fifoOut[35][10];
              muxOutConnector[36] = fifoOut[36][10];
              muxOutConnector[37] = fifoOut[37][10];
              muxOutConnector[38] = fifoOut[38][10];
              muxOutConnector[39] = fifoOut[39][10];
              muxOutConnector[40] = fifoOut[40][10];
              muxOutConnector[41] = fifoOut[41][10];
              muxOutConnector[42] = fifoOut[42][10];
              muxOutConnector[43] = fifoOut[43][10];
              muxOutConnector[44] = fifoOut[44][10];
              muxOutConnector[45] = fifoOut[45][10];
              muxOutConnector[46] = fifoOut[46][10];
              muxOutConnector[47] = fifoOut[47][10];
              muxOutConnector[48] = fifoOut[48][10];
              muxOutConnector[49] = fifoOut[49][10];
              muxOutConnector[50] = fifoOut[50][10];
              muxOutConnector[51] = fifoOut[51][10];
       end
       3: begin
              muxOutConnector[0] = fifoOut[38][4];
              muxOutConnector[1] = fifoOut[39][4];
              muxOutConnector[2] = fifoOut[40][4];
              muxOutConnector[3] = fifoOut[41][4];
              muxOutConnector[4] = fifoOut[42][4];
              muxOutConnector[5] = fifoOut[43][4];
              muxOutConnector[6] = fifoOut[44][4];
              muxOutConnector[7] = fifoOut[45][4];
              muxOutConnector[8] = fifoOut[46][4];
              muxOutConnector[9] = fifoOut[47][4];
              muxOutConnector[10] = fifoOut[48][4];
              muxOutConnector[11] = fifoOut[49][4];
              muxOutConnector[12] = fifoOut[50][4];
              muxOutConnector[13] = fifoOut[51][4];
              muxOutConnector[14] = fifoOut[26][3];
              muxOutConnector[15] = fifoOut[27][3];
              muxOutConnector[16] = fifoOut[28][3];
              muxOutConnector[17] = fifoOut[29][3];
              muxOutConnector[18] = fifoOut[30][3];
              muxOutConnector[19] = fifoOut[31][3];
              muxOutConnector[20] = fifoOut[32][3];
              muxOutConnector[21] = fifoOut[33][3];
              muxOutConnector[22] = fifoOut[34][3];
              muxOutConnector[23] = fifoOut[35][3];
              muxOutConnector[24] = fifoOut[36][3];
              muxOutConnector[25] = fifoOut[37][3];
              muxOutConnector[26] = fifoOut[26][10];
              muxOutConnector[27] = fifoOut[27][10];
              muxOutConnector[28] = fifoOut[28][10];
              muxOutConnector[29] = fifoOut[29][10];
              muxOutConnector[30] = fifoOut[30][10];
              muxOutConnector[31] = fifoOut[31][10];
              muxOutConnector[32] = fifoOut[32][10];
              muxOutConnector[33] = fifoOut[33][10];
              muxOutConnector[34] = fifoOut[34][10];
              muxOutConnector[35] = fifoOut[35][10];
              muxOutConnector[36] = fifoOut[36][10];
              muxOutConnector[37] = fifoOut[37][10];
              muxOutConnector[38] = fifoOut[38][10];
              muxOutConnector[39] = fifoOut[39][10];
              muxOutConnector[40] = fifoOut[40][10];
              muxOutConnector[41] = fifoOut[41][10];
              muxOutConnector[42] = fifoOut[42][10];
              muxOutConnector[43] = fifoOut[43][10];
              muxOutConnector[44] = fifoOut[44][10];
              muxOutConnector[45] = fifoOut[45][10];
              muxOutConnector[46] = fifoOut[46][10];
              muxOutConnector[47] = fifoOut[47][10];
              muxOutConnector[48] = fifoOut[48][10];
              muxOutConnector[49] = fifoOut[49][10];
              muxOutConnector[50] = fifoOut[50][10];
              muxOutConnector[51] = fifoOut[51][10];
       end
       4: begin
              muxOutConnector[0] = fifoOut[38][4];
              muxOutConnector[1] = fifoOut[39][4];
              muxOutConnector[2] = fifoOut[40][4];
              muxOutConnector[3] = fifoOut[41][4];
              muxOutConnector[4] = fifoOut[42][4];
              muxOutConnector[5] = fifoOut[19][3];
              muxOutConnector[6] = fifoOut[20][3];
              muxOutConnector[7] = fifoOut[21][3];
              muxOutConnector[8] = fifoOut[22][3];
              muxOutConnector[9] = fifoOut[23][3];
              muxOutConnector[10] = fifoOut[24][3];
              muxOutConnector[11] = fifoOut[25][3];
              muxOutConnector[12] = fifoOut[0][2];
              muxOutConnector[13] = fifoOut[1][2];
              muxOutConnector[14] = fifoOut[2][2];
              muxOutConnector[15] = fifoOut[3][2];
              muxOutConnector[16] = fifoOut[4][2];
              muxOutConnector[17] = fifoOut[5][2];
              muxOutConnector[18] = fifoOut[6][2];
              muxOutConnector[19] = fifoOut[7][2];
              muxOutConnector[20] = fifoOut[8][2];
              muxOutConnector[21] = fifoOut[9][2];
              muxOutConnector[22] = fifoOut[10][2];
              muxOutConnector[23] = fifoOut[11][2];
              muxOutConnector[24] = fifoOut[12][2];
              muxOutConnector[25] = fifoOut[13][2];
              muxOutConnector[26] = fifoOut[26][10];
              muxOutConnector[27] = fifoOut[27][10];
              muxOutConnector[28] = fifoOut[28][10];
              muxOutConnector[29] = fifoOut[29][10];
              muxOutConnector[30] = fifoOut[30][10];
              muxOutConnector[31] = fifoOut[31][10];
              muxOutConnector[32] = fifoOut[32][10];
              muxOutConnector[33] = fifoOut[33][10];
              muxOutConnector[34] = fifoOut[34][10];
              muxOutConnector[35] = fifoOut[35][10];
              muxOutConnector[36] = fifoOut[36][10];
              muxOutConnector[37] = fifoOut[37][10];
              muxOutConnector[38] = fifoOut[38][10];
              muxOutConnector[39] = fifoOut[39][10];
              muxOutConnector[40] = fifoOut[40][10];
              muxOutConnector[41] = fifoOut[41][10];
              muxOutConnector[42] = fifoOut[42][10];
              muxOutConnector[43] = fifoOut[43][10];
              muxOutConnector[44] = fifoOut[44][10];
              muxOutConnector[45] = fifoOut[45][10];
              muxOutConnector[46] = fifoOut[46][10];
              muxOutConnector[47] = fifoOut[47][10];
              muxOutConnector[48] = fifoOut[48][10];
              muxOutConnector[49] = fifoOut[49][10];
              muxOutConnector[50] = fifoOut[50][10];
              muxOutConnector[51] = fifoOut[51][10];
       end
       5: begin
              muxOutConnector[0] = fifoOut[14][3];
              muxOutConnector[1] = fifoOut[15][3];
              muxOutConnector[2] = fifoOut[16][3];
              muxOutConnector[3] = fifoOut[17][3];
              muxOutConnector[4] = fifoOut[18][3];
              muxOutConnector[5] = fifoOut[19][3];
              muxOutConnector[6] = fifoOut[20][3];
              muxOutConnector[7] = fifoOut[21][3];
              muxOutConnector[8] = fifoOut[22][3];
              muxOutConnector[9] = fifoOut[23][3];
              muxOutConnector[10] = fifoOut[24][3];
              muxOutConnector[11] = fifoOut[25][3];
              muxOutConnector[12] = fifoOut[0][2];
              muxOutConnector[13] = fifoOut[1][2];
              muxOutConnector[14] = fifoOut[2][2];
              muxOutConnector[15] = fifoOut[3][2];
              muxOutConnector[16] = fifoOut[4][2];
              muxOutConnector[17] = fifoOut[5][2];
              muxOutConnector[18] = fifoOut[6][2];
              muxOutConnector[19] = fifoOut[7][2];
              muxOutConnector[20] = fifoOut[8][2];
              muxOutConnector[21] = fifoOut[9][2];
              muxOutConnector[22] = fifoOut[10][2];
              muxOutConnector[23] = fifoOut[11][2];
              muxOutConnector[24] = fifoOut[12][2];
              muxOutConnector[25] = fifoOut[13][2];
              muxOutConnector[26] = fifoOut[26][10];
              muxOutConnector[27] = fifoOut[27][10];
              muxOutConnector[28] = fifoOut[28][10];
              muxOutConnector[29] = fifoOut[29][10];
              muxOutConnector[30] = fifoOut[30][10];
              muxOutConnector[31] = fifoOut[31][10];
              muxOutConnector[32] = fifoOut[32][10];
              muxOutConnector[33] = fifoOut[33][10];
              muxOutConnector[34] = fifoOut[34][10];
              muxOutConnector[35] = fifoOut[35][10];
              muxOutConnector[36] = fifoOut[36][10];
              muxOutConnector[37] = fifoOut[37][10];
              muxOutConnector[38] = fifoOut[38][10];
              muxOutConnector[39] = fifoOut[39][10];
              muxOutConnector[40] = fifoOut[40][10];
              muxOutConnector[41] = fifoOut[41][10];
              muxOutConnector[42] = fifoOut[42][10];
              muxOutConnector[43] = fifoOut[43][10];
              muxOutConnector[44] = fifoOut[44][10];
              muxOutConnector[45] = fifoOut[45][10];
              muxOutConnector[46] = fifoOut[46][10];
              muxOutConnector[47] = fifoOut[47][10];
              muxOutConnector[48] = fifoOut[48][10];
              muxOutConnector[49] = fifoOut[49][10];
              muxOutConnector[50] = fifoOut[50][10];
              muxOutConnector[51] = fifoOut[51][10];
       end
       6: begin
              muxOutConnector[0] = fifoOut[14][3];
              muxOutConnector[1] = fifoOut[15][3];
              muxOutConnector[2] = fifoOut[16][3];
              muxOutConnector[3] = fifoOut[17][3];
              muxOutConnector[4] = fifoOut[18][3];
              muxOutConnector[5] = fifoOut[19][3];
              muxOutConnector[6] = fifoOut[20][3];
              muxOutConnector[7] = fifoOut[21][3];
              muxOutConnector[8] = fifoOut[22][3];
              muxOutConnector[9] = fifoOut[23][3];
              muxOutConnector[10] = fifoOut[24][3];
              muxOutConnector[11] = fifoOut[25][3];
              muxOutConnector[12] = fifoOut[0][2];
              muxOutConnector[13] = fifoOut[1][2];
              muxOutConnector[14] = fifoOut[2][2];
              muxOutConnector[15] = fifoOut[3][2];
              muxOutConnector[16] = fifoOut[4][2];
              muxOutConnector[17] = fifoOut[5][2];
              muxOutConnector[18] = fifoOut[6][2];
              muxOutConnector[19] = fifoOut[7][2];
              muxOutConnector[20] = fifoOut[8][2];
              muxOutConnector[21] = fifoOut[9][2];
              muxOutConnector[22] = fifoOut[10][2];
              muxOutConnector[23] = fifoOut[11][2];
              muxOutConnector[24] = fifoOut[12][2];
              muxOutConnector[25] = fifoOut[13][2];
              muxOutConnector[26] = fifoOut[26][10];
              muxOutConnector[27] = fifoOut[27][10];
              muxOutConnector[28] = fifoOut[28][10];
              muxOutConnector[29] = fifoOut[29][10];
              muxOutConnector[30] = fifoOut[30][10];
              muxOutConnector[31] = fifoOut[31][10];
              muxOutConnector[32] = fifoOut[32][10];
              muxOutConnector[33] = fifoOut[33][10];
              muxOutConnector[34] = fifoOut[34][10];
              muxOutConnector[35] = fifoOut[35][10];
              muxOutConnector[36] = fifoOut[36][10];
              muxOutConnector[37] = fifoOut[37][10];
              muxOutConnector[38] = fifoOut[38][10];
              muxOutConnector[39] = fifoOut[39][10];
              muxOutConnector[40] = fifoOut[40][10];
              muxOutConnector[41] = fifoOut[41][10];
              muxOutConnector[42] = fifoOut[42][10];
              muxOutConnector[43] = fifoOut[43][10];
              muxOutConnector[44] = fifoOut[44][10];
              muxOutConnector[45] = fifoOut[45][10];
              muxOutConnector[46] = fifoOut[46][10];
              muxOutConnector[47] = fifoOut[47][10];
              muxOutConnector[48] = fifoOut[48][10];
              muxOutConnector[49] = fifoOut[49][10];
              muxOutConnector[50] = fifoOut[50][10];
              muxOutConnector[51] = fifoOut[51][10];
       end
       7: begin
              muxOutConnector[0] = fifoOut[14][3];
              muxOutConnector[1] = fifoOut[15][3];
              muxOutConnector[2] = fifoOut[16][3];
              muxOutConnector[3] = fifoOut[17][3];
              muxOutConnector[4] = fifoOut[18][3];
              muxOutConnector[5] = fifoOut[19][3];
              muxOutConnector[6] = fifoOut[20][3];
              muxOutConnector[7] = fifoOut[21][3];
              muxOutConnector[8] = fifoOut[22][3];
              muxOutConnector[9] = fifoOut[23][3];
              muxOutConnector[10] = fifoOut[24][3];
              muxOutConnector[11] = fifoOut[25][3];
              muxOutConnector[12] = fifoOut[0][2];
              muxOutConnector[13] = fifoOut[1][2];
              muxOutConnector[14] = fifoOut[2][2];
              muxOutConnector[15] = fifoOut[3][2];
              muxOutConnector[16] = fifoOut[4][2];
              muxOutConnector[17] = fifoOut[5][2];
              muxOutConnector[18] = fifoOut[6][2];
              muxOutConnector[19] = fifoOut[7][2];
              muxOutConnector[20] = fifoOut[8][2];
              muxOutConnector[21] = fifoOut[9][2];
              muxOutConnector[22] = fifoOut[10][2];
              muxOutConnector[23] = fifoOut[11][2];
              muxOutConnector[24] = fifoOut[12][2];
              muxOutConnector[25] = fifoOut[13][2];
              muxOutConnector[26] = fifoOut[26][10];
              muxOutConnector[27] = fifoOut[27][10];
              muxOutConnector[28] = fifoOut[28][10];
              muxOutConnector[29] = fifoOut[29][10];
              muxOutConnector[30] = fifoOut[30][10];
              muxOutConnector[31] = fifoOut[31][10];
              muxOutConnector[32] = fifoOut[32][10];
              muxOutConnector[33] = fifoOut[33][10];
              muxOutConnector[34] = fifoOut[34][10];
              muxOutConnector[35] = fifoOut[35][10];
              muxOutConnector[36] = fifoOut[36][10];
              muxOutConnector[37] = fifoOut[37][10];
              muxOutConnector[38] = fifoOut[38][10];
              muxOutConnector[39] = fifoOut[39][10];
              muxOutConnector[40] = fifoOut[40][10];
              muxOutConnector[41] = fifoOut[41][10];
              muxOutConnector[42] = fifoOut[42][10];
              muxOutConnector[43] = fifoOut[43][10];
              muxOutConnector[44] = fifoOut[44][10];
              muxOutConnector[45] = fifoOut[45][10];
              muxOutConnector[46] = fifoOut[46][10];
              muxOutConnector[47] = fifoOut[47][10];
              muxOutConnector[48] = fifoOut[48][10];
              muxOutConnector[49] = fifoOut[49][10];
              muxOutConnector[50] = fifoOut[50][10];
              muxOutConnector[51] = fifoOut[51][10];
       end
       8: begin
              muxOutConnector[0] = fifoOut[14][3];
              muxOutConnector[1] = fifoOut[15][3];
              muxOutConnector[2] = fifoOut[16][3];
              muxOutConnector[3] = fifoOut[17][3];
              muxOutConnector[4] = fifoOut[18][3];
              muxOutConnector[5] = fifoOut[19][3];
              muxOutConnector[6] = fifoOut[20][3];
              muxOutConnector[7] = fifoOut[21][3];
              muxOutConnector[8] = fifoOut[22][3];
              muxOutConnector[9] = fifoOut[23][3];
              muxOutConnector[10] = fifoOut[24][3];
              muxOutConnector[11] = fifoOut[25][3];
              muxOutConnector[12] = fifoOut[0][2];
              muxOutConnector[13] = fifoOut[1][2];
              muxOutConnector[14] = fifoOut[2][2];
              muxOutConnector[15] = fifoOut[3][2];
              muxOutConnector[16] = fifoOut[4][2];
              muxOutConnector[17] = fifoOut[5][2];
              muxOutConnector[18] = fifoOut[6][2];
              muxOutConnector[19] = fifoOut[7][2];
              muxOutConnector[20] = fifoOut[8][2];
              muxOutConnector[21] = fifoOut[9][2];
              muxOutConnector[22] = fifoOut[10][2];
              muxOutConnector[23] = fifoOut[11][2];
              muxOutConnector[24] = fifoOut[12][2];
              muxOutConnector[25] = fifoOut[13][2];
              muxOutConnector[26] = fifoOut[26][10];
              muxOutConnector[27] = fifoOut[27][10];
              muxOutConnector[28] = fifoOut[28][10];
              muxOutConnector[29] = fifoOut[29][10];
              muxOutConnector[30] = fifoOut[30][10];
              muxOutConnector[31] = fifoOut[31][10];
              muxOutConnector[32] = fifoOut[32][10];
              muxOutConnector[33] = fifoOut[33][10];
              muxOutConnector[34] = fifoOut[34][10];
              muxOutConnector[35] = fifoOut[35][10];
              muxOutConnector[36] = fifoOut[36][10];
              muxOutConnector[37] = fifoOut[37][10];
              muxOutConnector[38] = fifoOut[38][10];
              muxOutConnector[39] = fifoOut[39][10];
              muxOutConnector[40] = fifoOut[40][10];
              muxOutConnector[41] = fifoOut[41][10];
              muxOutConnector[42] = fifoOut[42][10];
              muxOutConnector[43] = fifoOut[43][10];
              muxOutConnector[44] = fifoOut[44][10];
              muxOutConnector[45] = fifoOut[45][10];
              muxOutConnector[46] = fifoOut[46][10];
              muxOutConnector[47] = fifoOut[47][10];
              muxOutConnector[48] = fifoOut[48][10];
              muxOutConnector[49] = fifoOut[49][10];
              muxOutConnector[50] = fifoOut[50][10];
              muxOutConnector[51] = fifoOut[51][10];
       end
       9: begin
              muxOutConnector[0] = fifoOut[14][3];
              muxOutConnector[1] = fifoOut[15][3];
              muxOutConnector[2] = fifoOut[16][3];
              muxOutConnector[3] = fifoOut[17][3];
              muxOutConnector[4] = fifoOut[18][3];
              muxOutConnector[5] = fifoOut[19][3];
              muxOutConnector[6] = fifoOut[20][3];
              muxOutConnector[7] = fifoOut[21][3];
              muxOutConnector[8] = fifoOut[22][3];
              muxOutConnector[9] = fifoOut[23][3];
              muxOutConnector[10] = fifoOut[24][3];
              muxOutConnector[11] = fifoOut[25][3];
              muxOutConnector[12] = fifoOut[0][2];
              muxOutConnector[13] = fifoOut[1][2];
              muxOutConnector[14] = fifoOut[2][2];
              muxOutConnector[15] = fifoOut[3][2];
              muxOutConnector[16] = fifoOut[4][2];
              muxOutConnector[17] = fifoOut[5][2];
              muxOutConnector[18] = fifoOut[6][2];
              muxOutConnector[19] = fifoOut[7][2];
              muxOutConnector[20] = fifoOut[8][2];
              muxOutConnector[21] = fifoOut[9][2];
              muxOutConnector[22] = fifoOut[10][2];
              muxOutConnector[23] = fifoOut[11][2];
              muxOutConnector[24] = fifoOut[12][2];
              muxOutConnector[25] = fifoOut[13][2];
              muxOutConnector[26] = fifoOut[26][10];
              muxOutConnector[27] = fifoOut[27][10];
              muxOutConnector[28] = fifoOut[28][10];
              muxOutConnector[29] = fifoOut[29][10];
              muxOutConnector[30] = fifoOut[30][10];
              muxOutConnector[31] = fifoOut[31][10];
              muxOutConnector[32] = fifoOut[32][10];
              muxOutConnector[33] = fifoOut[33][10];
              muxOutConnector[34] = fifoOut[34][10];
              muxOutConnector[35] = fifoOut[35][10];
              muxOutConnector[36] = fifoOut[36][10];
              muxOutConnector[37] = fifoOut[37][10];
              muxOutConnector[38] = fifoOut[38][10];
              muxOutConnector[39] = fifoOut[39][10];
              muxOutConnector[40] = fifoOut[40][10];
              muxOutConnector[41] = fifoOut[41][10];
              muxOutConnector[42] = fifoOut[42][10];
              muxOutConnector[43] = fifoOut[43][10];
              muxOutConnector[44] = fifoOut[44][10];
              muxOutConnector[45] = fifoOut[45][10];
              muxOutConnector[46] = fifoOut[46][10];
              muxOutConnector[47] = fifoOut[47][10];
              muxOutConnector[48] = fifoOut[48][10];
              muxOutConnector[49] = fifoOut[49][10];
              muxOutConnector[50] = fifoOut[50][10];
              muxOutConnector[51] = fifoOut[51][10];
       end
       10: begin
              muxOutConnector[0] = fifoOut[14][3];
              muxOutConnector[1] = fifoOut[15][3];
              muxOutConnector[2] = fifoOut[16][3];
              muxOutConnector[3] = fifoOut[17][3];
              muxOutConnector[4] = fifoOut[18][3];
              muxOutConnector[5] = fifoOut[19][3];
              muxOutConnector[6] = fifoOut[20][3];
              muxOutConnector[7] = fifoOut[21][3];
              muxOutConnector[8] = fifoOut[22][3];
              muxOutConnector[9] = fifoOut[23][3];
              muxOutConnector[10] = fifoOut[24][3];
              muxOutConnector[11] = fifoOut[25][3];
              muxOutConnector[12] = fifoOut[0][2];
              muxOutConnector[13] = fifoOut[1][2];
              muxOutConnector[14] = fifoOut[2][2];
              muxOutConnector[15] = fifoOut[3][2];
              muxOutConnector[16] = fifoOut[4][2];
              muxOutConnector[17] = fifoOut[5][2];
              muxOutConnector[18] = fifoOut[6][2];
              muxOutConnector[19] = fifoOut[7][2];
              muxOutConnector[20] = fifoOut[8][2];
              muxOutConnector[21] = fifoOut[9][2];
              muxOutConnector[22] = fifoOut[10][2];
              muxOutConnector[23] = fifoOut[11][2];
              muxOutConnector[24] = fifoOut[12][2];
              muxOutConnector[25] = fifoOut[13][2];
              muxOutConnector[26] = fifoOut[26][10];
              muxOutConnector[27] = fifoOut[27][10];
              muxOutConnector[28] = fifoOut[28][10];
              muxOutConnector[29] = fifoOut[29][10];
              muxOutConnector[30] = fifoOut[30][10];
              muxOutConnector[31] = fifoOut[31][10];
              muxOutConnector[32] = fifoOut[32][10];
              muxOutConnector[33] = fifoOut[33][10];
              muxOutConnector[34] = fifoOut[34][10];
              muxOutConnector[35] = fifoOut[35][10];
              muxOutConnector[36] = fifoOut[36][10];
              muxOutConnector[37] = fifoOut[37][10];
              muxOutConnector[38] = fifoOut[38][10];
              muxOutConnector[39] = fifoOut[39][10];
              muxOutConnector[40] = fifoOut[40][10];
              muxOutConnector[41] = fifoOut[41][10];
              muxOutConnector[42] = fifoOut[42][10];
              muxOutConnector[43] = fifoOut[19][9];
              muxOutConnector[44] = fifoOut[20][9];
              muxOutConnector[45] = fifoOut[21][9];
              muxOutConnector[46] = fifoOut[22][9];
              muxOutConnector[47] = fifoOut[23][9];
              muxOutConnector[48] = fifoOut[24][9];
              muxOutConnector[49] = fifoOut[25][9];
              muxOutConnector[50] = fifoOut[0][8];
              muxOutConnector[51] = fifoOut[1][8];
       end
       11: begin
              muxOutConnector[0] = fifoOut[14][3];
              muxOutConnector[1] = fifoOut[15][3];
              muxOutConnector[2] = fifoOut[16][3];
              muxOutConnector[3] = fifoOut[17][3];
              muxOutConnector[4] = fifoOut[18][3];
              muxOutConnector[5] = fifoOut[19][3];
              muxOutConnector[6] = fifoOut[20][3];
              muxOutConnector[7] = fifoOut[21][3];
              muxOutConnector[8] = fifoOut[22][3];
              muxOutConnector[9] = fifoOut[23][3];
              muxOutConnector[10] = fifoOut[24][3];
              muxOutConnector[11] = fifoOut[25][3];
              muxOutConnector[12] = fifoOut[0][2];
              muxOutConnector[13] = fifoOut[1][2];
              muxOutConnector[14] = fifoOut[2][2];
              muxOutConnector[15] = fifoOut[3][2];
              muxOutConnector[16] = fifoOut[4][2];
              muxOutConnector[17] = fifoOut[5][2];
              muxOutConnector[18] = fifoOut[6][2];
              muxOutConnector[19] = fifoOut[7][2];
              muxOutConnector[20] = fifoOut[8][2];
              muxOutConnector[21] = fifoOut[9][2];
              muxOutConnector[22] = fifoOut[10][2];
              muxOutConnector[23] = fifoOut[11][2];
              muxOutConnector[24] = fifoOut[12][2];
              muxOutConnector[25] = fifoOut[13][2];
              muxOutConnector[26] = fifoOut[2][9];
              muxOutConnector[27] = fifoOut[3][9];
              muxOutConnector[28] = fifoOut[4][9];
              muxOutConnector[29] = fifoOut[5][9];
              muxOutConnector[30] = fifoOut[6][9];
              muxOutConnector[31] = fifoOut[7][9];
              muxOutConnector[32] = fifoOut[8][9];
              muxOutConnector[33] = fifoOut[9][9];
              muxOutConnector[34] = fifoOut[10][9];
              muxOutConnector[35] = fifoOut[11][9];
              muxOutConnector[36] = fifoOut[12][9];
              muxOutConnector[37] = fifoOut[13][9];
              muxOutConnector[38] = fifoOut[14][9];
              muxOutConnector[39] = fifoOut[15][9];
              muxOutConnector[40] = fifoOut[16][9];
              muxOutConnector[41] = fifoOut[17][9];
              muxOutConnector[42] = fifoOut[18][9];
              muxOutConnector[43] = fifoOut[19][9];
              muxOutConnector[44] = fifoOut[20][9];
              muxOutConnector[45] = fifoOut[21][9];
              muxOutConnector[46] = fifoOut[22][9];
              muxOutConnector[47] = fifoOut[23][9];
              muxOutConnector[48] = fifoOut[24][9];
              muxOutConnector[49] = fifoOut[25][9];
              muxOutConnector[50] = fifoOut[0][8];
              muxOutConnector[51] = fifoOut[1][8];
       end
       12: begin
              muxOutConnector[0] = fifoOut[14][3];
              muxOutConnector[1] = fifoOut[15][3];
              muxOutConnector[2] = fifoOut[16][3];
              muxOutConnector[3] = fifoOut[17][3];
              muxOutConnector[4] = fifoOut[18][3];
              muxOutConnector[5] = fifoOut[26][11];
              muxOutConnector[6] = fifoOut[27][11];
              muxOutConnector[7] = fifoOut[28][11];
              muxOutConnector[8] = fifoOut[29][11];
              muxOutConnector[9] = fifoOut[30][11];
              muxOutConnector[10] = fifoOut[31][11];
              muxOutConnector[11] = fifoOut[32][11];
              muxOutConnector[12] = fifoOut[33][11];
              muxOutConnector[13] = fifoOut[34][11];
              muxOutConnector[14] = fifoOut[35][11];
              muxOutConnector[15] = fifoOut[36][11];
              muxOutConnector[16] = fifoOut[37][11];
              muxOutConnector[17] = fifoOut[38][11];
              muxOutConnector[18] = fifoOut[39][11];
              muxOutConnector[19] = fifoOut[40][11];
              muxOutConnector[20] = fifoOut[41][11];
              muxOutConnector[21] = fifoOut[42][11];
              muxOutConnector[22] = fifoOut[43][11];
              muxOutConnector[23] = fifoOut[44][11];
              muxOutConnector[24] = fifoOut[45][11];
              muxOutConnector[25] = fifoOut[46][11];
              muxOutConnector[26] = fifoOut[2][9];
              muxOutConnector[27] = fifoOut[3][9];
              muxOutConnector[28] = fifoOut[4][9];
              muxOutConnector[29] = fifoOut[5][9];
              muxOutConnector[30] = fifoOut[6][9];
              muxOutConnector[31] = fifoOut[7][9];
              muxOutConnector[32] = fifoOut[8][9];
              muxOutConnector[33] = fifoOut[9][9];
              muxOutConnector[34] = fifoOut[10][9];
              muxOutConnector[35] = fifoOut[11][9];
              muxOutConnector[36] = fifoOut[12][9];
              muxOutConnector[37] = fifoOut[13][9];
              muxOutConnector[38] = fifoOut[14][9];
              muxOutConnector[39] = fifoOut[15][9];
              muxOutConnector[40] = fifoOut[16][9];
              muxOutConnector[41] = fifoOut[17][9];
              muxOutConnector[42] = fifoOut[18][9];
              muxOutConnector[43] = fifoOut[19][9];
              muxOutConnector[44] = fifoOut[20][9];
              muxOutConnector[45] = fifoOut[21][9];
              muxOutConnector[46] = fifoOut[22][9];
              muxOutConnector[47] = fifoOut[23][9];
              muxOutConnector[48] = fifoOut[24][9];
              muxOutConnector[49] = fifoOut[25][9];
              muxOutConnector[50] = fifoOut[0][8];
              muxOutConnector[51] = fifoOut[1][8];
       end
       13: begin
              muxOutConnector[0] = fifoOut[14][3];
              muxOutConnector[1] = fifoOut[15][3];
              muxOutConnector[2] = fifoOut[16][3];
              muxOutConnector[3] = fifoOut[17][3];
              muxOutConnector[4] = fifoOut[18][3];
              muxOutConnector[5] = fifoOut[26][11];
              muxOutConnector[6] = fifoOut[27][11];
              muxOutConnector[7] = fifoOut[28][11];
              muxOutConnector[8] = fifoOut[29][11];
              muxOutConnector[9] = fifoOut[30][11];
              muxOutConnector[10] = fifoOut[31][11];
              muxOutConnector[11] = fifoOut[32][11];
              muxOutConnector[12] = fifoOut[33][11];
              muxOutConnector[13] = fifoOut[34][11];
              muxOutConnector[14] = fifoOut[35][11];
              muxOutConnector[15] = fifoOut[36][11];
              muxOutConnector[16] = fifoOut[37][11];
              muxOutConnector[17] = fifoOut[38][11];
              muxOutConnector[18] = fifoOut[39][11];
              muxOutConnector[19] = fifoOut[40][11];
              muxOutConnector[20] = fifoOut[41][11];
              muxOutConnector[21] = fifoOut[42][11];
              muxOutConnector[22] = fifoOut[43][11];
              muxOutConnector[23] = fifoOut[44][11];
              muxOutConnector[24] = fifoOut[45][11];
              muxOutConnector[25] = fifoOut[46][11];
              muxOutConnector[26] = fifoOut[2][9];
              muxOutConnector[27] = fifoOut[3][9];
              muxOutConnector[28] = fifoOut[4][9];
              muxOutConnector[29] = fifoOut[5][9];
              muxOutConnector[30] = fifoOut[6][9];
              muxOutConnector[31] = fifoOut[7][9];
              muxOutConnector[32] = fifoOut[8][9];
              muxOutConnector[33] = fifoOut[9][9];
              muxOutConnector[34] = fifoOut[10][9];
              muxOutConnector[35] = fifoOut[11][9];
              muxOutConnector[36] = fifoOut[12][9];
              muxOutConnector[37] = fifoOut[13][9];
              muxOutConnector[38] = fifoOut[14][9];
              muxOutConnector[39] = fifoOut[15][9];
              muxOutConnector[40] = fifoOut[16][9];
              muxOutConnector[41] = fifoOut[17][9];
              muxOutConnector[42] = fifoOut[18][9];
              muxOutConnector[43] = fifoOut[19][9];
              muxOutConnector[44] = fifoOut[20][9];
              muxOutConnector[45] = fifoOut[21][9];
              muxOutConnector[46] = fifoOut[22][9];
              muxOutConnector[47] = fifoOut[23][9];
              muxOutConnector[48] = fifoOut[24][9];
              muxOutConnector[49] = fifoOut[25][9];
              muxOutConnector[50] = fifoOut[0][8];
              muxOutConnector[51] = fifoOut[1][8];
       end
       14: begin
              muxOutConnector[0] = fifoOut[14][3];
              muxOutConnector[1] = fifoOut[15][3];
              muxOutConnector[2] = fifoOut[16][3];
              muxOutConnector[3] = fifoOut[17][3];
              muxOutConnector[4] = fifoOut[18][3];
              muxOutConnector[5] = fifoOut[26][11];
              muxOutConnector[6] = fifoOut[27][11];
              muxOutConnector[7] = fifoOut[28][11];
              muxOutConnector[8] = fifoOut[29][11];
              muxOutConnector[9] = fifoOut[30][11];
              muxOutConnector[10] = fifoOut[31][11];
              muxOutConnector[11] = fifoOut[32][11];
              muxOutConnector[12] = fifoOut[33][11];
              muxOutConnector[13] = fifoOut[34][11];
              muxOutConnector[14] = fifoOut[35][11];
              muxOutConnector[15] = fifoOut[36][11];
              muxOutConnector[16] = fifoOut[37][11];
              muxOutConnector[17] = fifoOut[38][11];
              muxOutConnector[18] = fifoOut[39][11];
              muxOutConnector[19] = fifoOut[40][11];
              muxOutConnector[20] = fifoOut[41][11];
              muxOutConnector[21] = fifoOut[42][11];
              muxOutConnector[22] = fifoOut[43][11];
              muxOutConnector[23] = fifoOut[44][11];
              muxOutConnector[24] = fifoOut[45][11];
              muxOutConnector[25] = fifoOut[46][11];
              muxOutConnector[26] = fifoOut[2][9];
              muxOutConnector[27] = fifoOut[3][9];
              muxOutConnector[28] = fifoOut[4][9];
              muxOutConnector[29] = fifoOut[5][9];
              muxOutConnector[30] = fifoOut[6][9];
              muxOutConnector[31] = fifoOut[7][9];
              muxOutConnector[32] = fifoOut[8][9];
              muxOutConnector[33] = fifoOut[9][9];
              muxOutConnector[34] = fifoOut[10][9];
              muxOutConnector[35] = fifoOut[11][9];
              muxOutConnector[36] = fifoOut[12][9];
              muxOutConnector[37] = fifoOut[13][9];
              muxOutConnector[38] = fifoOut[14][9];
              muxOutConnector[39] = fifoOut[15][9];
              muxOutConnector[40] = fifoOut[16][9];
              muxOutConnector[41] = fifoOut[17][9];
              muxOutConnector[42] = fifoOut[18][9];
              muxOutConnector[43] = fifoOut[19][9];
              muxOutConnector[44] = fifoOut[20][9];
              muxOutConnector[45] = fifoOut[21][9];
              muxOutConnector[46] = fifoOut[22][9];
              muxOutConnector[47] = fifoOut[23][9];
              muxOutConnector[48] = fifoOut[24][9];
              muxOutConnector[49] = fifoOut[25][9];
              muxOutConnector[50] = fifoOut[0][8];
              muxOutConnector[51] = fifoOut[1][8];
       end
       15: begin
              muxOutConnector[0] = fifoOut[14][3];
              muxOutConnector[1] = fifoOut[15][3];
              muxOutConnector[2] = fifoOut[16][3];
              muxOutConnector[3] = fifoOut[50][0];
              muxOutConnector[4] = fifoOut[51][0];
              muxOutConnector[5] = fifoOut[26][11];
              muxOutConnector[6] = fifoOut[27][11];
              muxOutConnector[7] = fifoOut[28][11];
              muxOutConnector[8] = fifoOut[29][11];
              muxOutConnector[9] = fifoOut[30][11];
              muxOutConnector[10] = fifoOut[31][11];
              muxOutConnector[11] = fifoOut[32][11];
              muxOutConnector[12] = fifoOut[33][11];
              muxOutConnector[13] = fifoOut[34][11];
              muxOutConnector[14] = fifoOut[35][11];
              muxOutConnector[15] = fifoOut[36][11];
              muxOutConnector[16] = fifoOut[37][11];
              muxOutConnector[17] = fifoOut[38][11];
              muxOutConnector[18] = fifoOut[39][11];
              muxOutConnector[19] = fifoOut[40][11];
              muxOutConnector[20] = fifoOut[41][11];
              muxOutConnector[21] = fifoOut[42][11];
              muxOutConnector[22] = fifoOut[43][11];
              muxOutConnector[23] = fifoOut[44][11];
              muxOutConnector[24] = fifoOut[45][11];
              muxOutConnector[25] = fifoOut[46][11];
              muxOutConnector[26] = fifoOut[2][9];
              muxOutConnector[27] = fifoOut[3][9];
              muxOutConnector[28] = fifoOut[4][9];
              muxOutConnector[29] = fifoOut[5][9];
              muxOutConnector[30] = fifoOut[6][9];
              muxOutConnector[31] = fifoOut[7][9];
              muxOutConnector[32] = fifoOut[8][9];
              muxOutConnector[33] = fifoOut[9][9];
              muxOutConnector[34] = fifoOut[10][9];
              muxOutConnector[35] = fifoOut[11][9];
              muxOutConnector[36] = fifoOut[12][9];
              muxOutConnector[37] = fifoOut[13][9];
              muxOutConnector[38] = fifoOut[14][9];
              muxOutConnector[39] = fifoOut[15][9];
              muxOutConnector[40] = fifoOut[16][9];
              muxOutConnector[41] = fifoOut[17][9];
              muxOutConnector[42] = fifoOut[18][9];
              muxOutConnector[43] = fifoOut[19][9];
              muxOutConnector[44] = fifoOut[20][9];
              muxOutConnector[45] = fifoOut[21][9];
              muxOutConnector[46] = fifoOut[22][9];
              muxOutConnector[47] = fifoOut[23][9];
              muxOutConnector[48] = fifoOut[24][9];
              muxOutConnector[49] = fifoOut[25][9];
              muxOutConnector[50] = fifoOut[0][8];
              muxOutConnector[51] = fifoOut[1][8];
       end
       16: begin
              muxOutConnector[0] = fifoOut[47][0];
              muxOutConnector[1] = fifoOut[48][0];
              muxOutConnector[2] = fifoOut[49][0];
              muxOutConnector[3] = fifoOut[50][0];
              muxOutConnector[4] = fifoOut[51][0];
              muxOutConnector[5] = fifoOut[26][11];
              muxOutConnector[6] = fifoOut[27][11];
              muxOutConnector[7] = fifoOut[28][11];
              muxOutConnector[8] = fifoOut[29][11];
              muxOutConnector[9] = fifoOut[30][11];
              muxOutConnector[10] = fifoOut[31][11];
              muxOutConnector[11] = fifoOut[32][11];
              muxOutConnector[12] = fifoOut[33][11];
              muxOutConnector[13] = fifoOut[34][11];
              muxOutConnector[14] = fifoOut[35][11];
              muxOutConnector[15] = fifoOut[36][11];
              muxOutConnector[16] = fifoOut[37][11];
              muxOutConnector[17] = fifoOut[38][11];
              muxOutConnector[18] = fifoOut[39][11];
              muxOutConnector[19] = fifoOut[40][11];
              muxOutConnector[20] = fifoOut[41][11];
              muxOutConnector[21] = fifoOut[42][11];
              muxOutConnector[22] = fifoOut[43][11];
              muxOutConnector[23] = fifoOut[44][11];
              muxOutConnector[24] = fifoOut[45][11];
              muxOutConnector[25] = fifoOut[46][11];
              muxOutConnector[26] = fifoOut[2][9];
              muxOutConnector[27] = fifoOut[3][9];
              muxOutConnector[28] = fifoOut[4][9];
              muxOutConnector[29] = fifoOut[5][9];
              muxOutConnector[30] = fifoOut[6][9];
              muxOutConnector[31] = fifoOut[7][9];
              muxOutConnector[32] = fifoOut[8][9];
              muxOutConnector[33] = fifoOut[9][9];
              muxOutConnector[34] = fifoOut[10][9];
              muxOutConnector[35] = fifoOut[11][9];
              muxOutConnector[36] = fifoOut[12][9];
              muxOutConnector[37] = fifoOut[13][9];
              muxOutConnector[38] = fifoOut[14][9];
              muxOutConnector[39] = fifoOut[15][9];
              muxOutConnector[40] = fifoOut[16][9];
              muxOutConnector[41] = fifoOut[17][9];
              muxOutConnector[42] = fifoOut[18][9];
              muxOutConnector[43] = fifoOut[19][9];
              muxOutConnector[44] = fifoOut[20][9];
              muxOutConnector[45] = fifoOut[21][9];
              muxOutConnector[46] = fifoOut[22][9];
              muxOutConnector[47] = fifoOut[23][9];
              muxOutConnector[48] = fifoOut[24][9];
              muxOutConnector[49] = fifoOut[25][9];
              muxOutConnector[50] = fifoOut[0][8];
              muxOutConnector[51] = fifoOut[1][8];
       end
       17: begin
              muxOutConnector[0] = fifoOut[47][0];
              muxOutConnector[1] = fifoOut[48][0];
              muxOutConnector[2] = fifoOut[49][0];
              muxOutConnector[3] = fifoOut[50][0];
              muxOutConnector[4] = fifoOut[51][0];
              muxOutConnector[5] = fifoOut[26][11];
              muxOutConnector[6] = fifoOut[27][11];
              muxOutConnector[7] = fifoOut[28][11];
              muxOutConnector[8] = fifoOut[29][11];
              muxOutConnector[9] = fifoOut[30][11];
              muxOutConnector[10] = fifoOut[31][11];
              muxOutConnector[11] = fifoOut[32][11];
              muxOutConnector[12] = fifoOut[33][11];
              muxOutConnector[13] = fifoOut[34][11];
              muxOutConnector[14] = fifoOut[35][11];
              muxOutConnector[15] = fifoOut[36][11];
              muxOutConnector[16] = fifoOut[37][11];
              muxOutConnector[17] = fifoOut[38][11];
              muxOutConnector[18] = fifoOut[39][11];
              muxOutConnector[19] = fifoOut[40][11];
              muxOutConnector[20] = fifoOut[41][11];
              muxOutConnector[21] = fifoOut[42][11];
              muxOutConnector[22] = fifoOut[43][11];
              muxOutConnector[23] = fifoOut[44][11];
              muxOutConnector[24] = fifoOut[45][11];
              muxOutConnector[25] = fifoOut[46][11];
              muxOutConnector[26] = fifoOut[2][9];
              muxOutConnector[27] = fifoOut[3][9];
              muxOutConnector[28] = fifoOut[4][9];
              muxOutConnector[29] = fifoOut[5][9];
              muxOutConnector[30] = fifoOut[6][9];
              muxOutConnector[31] = fifoOut[7][9];
              muxOutConnector[32] = fifoOut[8][9];
              muxOutConnector[33] = fifoOut[9][9];
              muxOutConnector[34] = fifoOut[10][9];
              muxOutConnector[35] = fifoOut[11][9];
              muxOutConnector[36] = fifoOut[12][9];
              muxOutConnector[37] = fifoOut[13][9];
              muxOutConnector[38] = fifoOut[14][9];
              muxOutConnector[39] = fifoOut[15][9];
              muxOutConnector[40] = fifoOut[16][9];
              muxOutConnector[41] = fifoOut[17][9];
              muxOutConnector[42] = fifoOut[18][9];
              muxOutConnector[43] = fifoOut[19][9];
              muxOutConnector[44] = fifoOut[20][9];
              muxOutConnector[45] = fifoOut[21][9];
              muxOutConnector[46] = fifoOut[22][9];
              muxOutConnector[47] = fifoOut[23][9];
              muxOutConnector[48] = fifoOut[24][9];
              muxOutConnector[49] = fifoOut[25][9];
              muxOutConnector[50] = fifoOut[0][8];
              muxOutConnector[51] = fifoOut[1][8];
       end
       18: begin
              muxOutConnector[0] = fifoOut[47][0];
              muxOutConnector[1] = fifoOut[48][0];
              muxOutConnector[2] = fifoOut[49][0];
              muxOutConnector[3] = fifoOut[50][0];
              muxOutConnector[4] = fifoOut[51][0];
              muxOutConnector[5] = fifoOut[26][11];
              muxOutConnector[6] = fifoOut[27][11];
              muxOutConnector[7] = fifoOut[28][11];
              muxOutConnector[8] = fifoOut[29][11];
              muxOutConnector[9] = fifoOut[30][11];
              muxOutConnector[10] = fifoOut[31][11];
              muxOutConnector[11] = fifoOut[32][11];
              muxOutConnector[12] = fifoOut[33][11];
              muxOutConnector[13] = fifoOut[34][11];
              muxOutConnector[14] = fifoOut[35][11];
              muxOutConnector[15] = fifoOut[36][11];
              muxOutConnector[16] = fifoOut[37][11];
              muxOutConnector[17] = fifoOut[38][11];
              muxOutConnector[18] = fifoOut[39][11];
              muxOutConnector[19] = fifoOut[40][11];
              muxOutConnector[20] = fifoOut[41][11];
              muxOutConnector[21] = fifoOut[42][11];
              muxOutConnector[22] = fifoOut[43][11];
              muxOutConnector[23] = fifoOut[44][11];
              muxOutConnector[24] = fifoOut[45][11];
              muxOutConnector[25] = fifoOut[46][11];
              muxOutConnector[26] = fifoOut[2][9];
              muxOutConnector[27] = fifoOut[3][9];
              muxOutConnector[28] = fifoOut[4][9];
              muxOutConnector[29] = fifoOut[5][9];
              muxOutConnector[30] = fifoOut[6][9];
              muxOutConnector[31] = fifoOut[7][9];
              muxOutConnector[32] = fifoOut[8][9];
              muxOutConnector[33] = fifoOut[9][9];
              muxOutConnector[34] = fifoOut[10][9];
              muxOutConnector[35] = fifoOut[11][9];
              muxOutConnector[36] = fifoOut[12][9];
              muxOutConnector[37] = fifoOut[13][9];
              muxOutConnector[38] = fifoOut[14][9];
              muxOutConnector[39] = fifoOut[15][9];
              muxOutConnector[40] = fifoOut[16][9];
              muxOutConnector[41] = fifoOut[17][9];
              muxOutConnector[42] = fifoOut[18][9];
              muxOutConnector[43] = fifoOut[19][9];
              muxOutConnector[44] = fifoOut[20][9];
              muxOutConnector[45] = fifoOut[21][9];
              muxOutConnector[46] = fifoOut[22][9];
              muxOutConnector[47] = fifoOut[23][9];
              muxOutConnector[48] = fifoOut[24][9];
              muxOutConnector[49] = fifoOut[25][9];
              muxOutConnector[50] = fifoOut[0][8];
              muxOutConnector[51] = fifoOut[1][8];
       end
       19: begin
              muxOutConnector[0] = fifoOut[47][0];
              muxOutConnector[1] = fifoOut[48][0];
              muxOutConnector[2] = fifoOut[49][0];
              muxOutConnector[3] = fifoOut[50][0];
              muxOutConnector[4] = fifoOut[51][0];
              muxOutConnector[5] = fifoOut[26][11];
              muxOutConnector[6] = fifoOut[27][11];
              muxOutConnector[7] = fifoOut[28][11];
              muxOutConnector[8] = fifoOut[29][11];
              muxOutConnector[9] = fifoOut[30][11];
              muxOutConnector[10] = fifoOut[31][11];
              muxOutConnector[11] = fifoOut[32][11];
              muxOutConnector[12] = fifoOut[33][11];
              muxOutConnector[13] = fifoOut[34][11];
              muxOutConnector[14] = fifoOut[35][11];
              muxOutConnector[15] = fifoOut[36][11];
              muxOutConnector[16] = fifoOut[37][11];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[2][9];
              muxOutConnector[27] = fifoOut[3][9];
              muxOutConnector[28] = fifoOut[4][9];
              muxOutConnector[29] = fifoOut[5][9];
              muxOutConnector[30] = fifoOut[6][9];
              muxOutConnector[31] = fifoOut[7][9];
              muxOutConnector[32] = fifoOut[8][9];
              muxOutConnector[33] = fifoOut[9][9];
              muxOutConnector[34] = fifoOut[10][9];
              muxOutConnector[35] = fifoOut[11][9];
              muxOutConnector[36] = fifoOut[12][9];
              muxOutConnector[37] = fifoOut[13][9];
              muxOutConnector[38] = fifoOut[14][9];
              muxOutConnector[39] = fifoOut[15][9];
              muxOutConnector[40] = fifoOut[16][9];
              muxOutConnector[41] = fifoOut[17][9];
              muxOutConnector[42] = fifoOut[18][9];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
