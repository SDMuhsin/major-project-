`timescale 1ns / 1ps
module LMem1To0_511_circ5_ys_yu_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        wr_en,
        feedback_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 13;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input [ADDRESSWIDTH-1:0]unloadAddress;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

input feedback_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        if(feedback_en) begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= fifoOut[i][c-1];
         end
        end
        else begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= ly0InConnector[i];
         end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
       0: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = fifoOut[21][11][w-1];
              unloadMuxOut[28] = fifoOut[22][11][w-1];
              unloadMuxOut[29] = fifoOut[23][11][w-1];
              unloadMuxOut[30] = fifoOut[24][11][w-1];
              unloadMuxOut[31] = fifoOut[25][11][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[0][10][w-1];
              unloadMuxOut[1] = fifoOut[1][10][w-1];
              unloadMuxOut[2] = fifoOut[2][10][w-1];
              unloadMuxOut[3] = fifoOut[3][10][w-1];
              unloadMuxOut[4] = fifoOut[4][10][w-1];
              unloadMuxOut[5] = fifoOut[5][10][w-1];
              unloadMuxOut[6] = fifoOut[6][10][w-1];
              unloadMuxOut[7] = fifoOut[7][10][w-1];
              unloadMuxOut[8] = fifoOut[8][10][w-1];
              unloadMuxOut[9] = fifoOut[9][10][w-1];
              unloadMuxOut[10] = fifoOut[10][10][w-1];
              unloadMuxOut[11] = fifoOut[11][10][w-1];
              unloadMuxOut[12] = fifoOut[12][10][w-1];
              unloadMuxOut[13] = fifoOut[13][10][w-1];
              unloadMuxOut[14] = fifoOut[14][10][w-1];
              unloadMuxOut[15] = fifoOut[15][10][w-1];
              unloadMuxOut[16] = fifoOut[16][10][w-1];
              unloadMuxOut[17] = fifoOut[17][10][w-1];
              unloadMuxOut[18] = fifoOut[18][10][w-1];
              unloadMuxOut[19] = fifoOut[19][10][w-1];
              unloadMuxOut[20] = fifoOut[20][10][w-1];
              unloadMuxOut[21] = fifoOut[21][10][w-1];
              unloadMuxOut[22] = fifoOut[22][10][w-1];
              unloadMuxOut[23] = fifoOut[23][10][w-1];
              unloadMuxOut[24] = fifoOut[24][10][w-1];
              unloadMuxOut[25] = fifoOut[25][10][w-1];
              unloadMuxOut[26] = fifoOut[0][9][w-1];
              unloadMuxOut[27] = fifoOut[1][9][w-1];
              unloadMuxOut[28] = fifoOut[2][9][w-1];
              unloadMuxOut[29] = fifoOut[3][9][w-1];
              unloadMuxOut[30] = fifoOut[4][9][w-1];
              unloadMuxOut[31] = fifoOut[5][9][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[6][9][w-1];
              unloadMuxOut[1] = fifoOut[7][9][w-1];
              unloadMuxOut[2] = fifoOut[8][9][w-1];
              unloadMuxOut[3] = fifoOut[9][9][w-1];
              unloadMuxOut[4] = fifoOut[10][9][w-1];
              unloadMuxOut[5] = fifoOut[11][9][w-1];
              unloadMuxOut[6] = fifoOut[12][9][w-1];
              unloadMuxOut[7] = fifoOut[13][9][w-1];
              unloadMuxOut[8] = fifoOut[14][9][w-1];
              unloadMuxOut[9] = fifoOut[15][9][w-1];
              unloadMuxOut[10] = fifoOut[16][9][w-1];
              unloadMuxOut[11] = fifoOut[17][9][w-1];
              unloadMuxOut[12] = fifoOut[18][9][w-1];
              unloadMuxOut[13] = fifoOut[19][9][w-1];
              unloadMuxOut[14] = fifoOut[20][9][w-1];
              unloadMuxOut[15] = fifoOut[21][9][w-1];
              unloadMuxOut[16] = fifoOut[22][9][w-1];
              unloadMuxOut[17] = fifoOut[23][9][w-1];
              unloadMuxOut[18] = fifoOut[24][9][w-1];
              unloadMuxOut[19] = fifoOut[25][9][w-1];
              unloadMuxOut[20] = fifoOut[0][8][w-1];
              unloadMuxOut[21] = fifoOut[1][8][w-1];
              unloadMuxOut[22] = fifoOut[2][8][w-1];
              unloadMuxOut[23] = fifoOut[3][8][w-1];
              unloadMuxOut[24] = fifoOut[4][8][w-1];
              unloadMuxOut[25] = fifoOut[5][8][w-1];
              unloadMuxOut[26] = fifoOut[6][8][w-1];
              unloadMuxOut[27] = fifoOut[7][8][w-1];
              unloadMuxOut[28] = fifoOut[8][8][w-1];
              unloadMuxOut[29] = fifoOut[9][8][w-1];
              unloadMuxOut[30] = fifoOut[10][8][w-1];
              unloadMuxOut[31] = fifoOut[11][8][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[12][8][w-1];
              unloadMuxOut[1] = fifoOut[13][8][w-1];
              unloadMuxOut[2] = fifoOut[14][8][w-1];
              unloadMuxOut[3] = fifoOut[15][8][w-1];
              unloadMuxOut[4] = fifoOut[16][8][w-1];
              unloadMuxOut[5] = fifoOut[17][8][w-1];
              unloadMuxOut[6] = fifoOut[18][8][w-1];
              unloadMuxOut[7] = fifoOut[19][8][w-1];
              unloadMuxOut[8] = fifoOut[20][8][w-1];
              unloadMuxOut[9] = fifoOut[21][8][w-1];
              unloadMuxOut[10] = fifoOut[22][8][w-1];
              unloadMuxOut[11] = fifoOut[23][8][w-1];
              unloadMuxOut[12] = fifoOut[24][8][w-1];
              unloadMuxOut[13] = fifoOut[25][8][w-1];
              unloadMuxOut[14] = fifoOut[0][7][w-1];
              unloadMuxOut[15] = fifoOut[1][7][w-1];
              unloadMuxOut[16] = fifoOut[2][7][w-1];
              unloadMuxOut[17] = fifoOut[3][7][w-1];
              unloadMuxOut[18] = fifoOut[4][7][w-1];
              unloadMuxOut[19] = fifoOut[5][7][w-1];
              unloadMuxOut[20] = fifoOut[6][7][w-1];
              unloadMuxOut[21] = fifoOut[7][7][w-1];
              unloadMuxOut[22] = fifoOut[8][7][w-1];
              unloadMuxOut[23] = fifoOut[9][7][w-1];
              unloadMuxOut[24] = fifoOut[10][7][w-1];
              unloadMuxOut[25] = fifoOut[11][7][w-1];
              unloadMuxOut[26] = fifoOut[12][7][w-1];
              unloadMuxOut[27] = fifoOut[13][7][w-1];
              unloadMuxOut[28] = fifoOut[14][7][w-1];
              unloadMuxOut[29] = fifoOut[15][7][w-1];
              unloadMuxOut[30] = fifoOut[16][7][w-1];
              unloadMuxOut[31] = fifoOut[17][7][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[18][7][w-1];
              unloadMuxOut[1] = fifoOut[19][7][w-1];
              unloadMuxOut[2] = fifoOut[20][7][w-1];
              unloadMuxOut[3] = fifoOut[21][7][w-1];
              unloadMuxOut[4] = fifoOut[22][7][w-1];
              unloadMuxOut[5] = fifoOut[23][7][w-1];
              unloadMuxOut[6] = fifoOut[24][7][w-1];
              unloadMuxOut[7] = fifoOut[25][7][w-1];
              unloadMuxOut[8] = fifoOut[0][6][w-1];
              unloadMuxOut[9] = fifoOut[1][6][w-1];
              unloadMuxOut[10] = fifoOut[2][6][w-1];
              unloadMuxOut[11] = fifoOut[3][6][w-1];
              unloadMuxOut[12] = fifoOut[4][6][w-1];
              unloadMuxOut[13] = fifoOut[5][6][w-1];
              unloadMuxOut[14] = fifoOut[6][6][w-1];
              unloadMuxOut[15] = fifoOut[7][6][w-1];
              unloadMuxOut[16] = fifoOut[8][6][w-1];
              unloadMuxOut[17] = fifoOut[9][6][w-1];
              unloadMuxOut[18] = fifoOut[10][6][w-1];
              unloadMuxOut[19] = fifoOut[11][6][w-1];
              unloadMuxOut[20] = fifoOut[12][6][w-1];
              unloadMuxOut[21] = fifoOut[13][6][w-1];
              unloadMuxOut[22] = fifoOut[14][6][w-1];
              unloadMuxOut[23] = fifoOut[15][6][w-1];
              unloadMuxOut[24] = fifoOut[16][6][w-1];
              unloadMuxOut[25] = fifoOut[17][6][w-1];
              unloadMuxOut[26] = fifoOut[18][6][w-1];
              unloadMuxOut[27] = fifoOut[19][6][w-1];
              unloadMuxOut[28] = fifoOut[20][6][w-1];
              unloadMuxOut[29] = fifoOut[21][6][w-1];
              unloadMuxOut[30] = fifoOut[22][6][w-1];
              unloadMuxOut[31] = fifoOut[23][6][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[24][6][w-1];
              unloadMuxOut[1] = fifoOut[25][6][w-1];
              unloadMuxOut[2] = fifoOut[0][5][w-1];
              unloadMuxOut[3] = fifoOut[1][5][w-1];
              unloadMuxOut[4] = fifoOut[2][5][w-1];
              unloadMuxOut[5] = fifoOut[3][5][w-1];
              unloadMuxOut[6] = fifoOut[4][5][w-1];
              unloadMuxOut[7] = fifoOut[5][5][w-1];
              unloadMuxOut[8] = fifoOut[6][5][w-1];
              unloadMuxOut[9] = fifoOut[7][5][w-1];
              unloadMuxOut[10] = fifoOut[8][5][w-1];
              unloadMuxOut[11] = fifoOut[9][5][w-1];
              unloadMuxOut[12] = fifoOut[10][5][w-1];
              unloadMuxOut[13] = fifoOut[11][5][w-1];
              unloadMuxOut[14] = fifoOut[12][5][w-1];
              unloadMuxOut[15] = fifoOut[13][5][w-1];
              unloadMuxOut[16] = fifoOut[14][5][w-1];
              unloadMuxOut[17] = fifoOut[15][5][w-1];
              unloadMuxOut[18] = fifoOut[16][5][w-1];
              unloadMuxOut[19] = fifoOut[26][12][w-1];
              unloadMuxOut[20] = fifoOut[27][12][w-1];
              unloadMuxOut[21] = fifoOut[28][12][w-1];
              unloadMuxOut[22] = fifoOut[29][12][w-1];
              unloadMuxOut[23] = fifoOut[30][12][w-1];
              unloadMuxOut[24] = fifoOut[31][12][w-1];
              unloadMuxOut[25] = fifoOut[32][12][w-1];
              unloadMuxOut[26] = fifoOut[33][12][w-1];
              unloadMuxOut[27] = fifoOut[34][12][w-1];
              unloadMuxOut[28] = fifoOut[35][12][w-1];
              unloadMuxOut[29] = fifoOut[36][12][w-1];
              unloadMuxOut[30] = fifoOut[37][12][w-1];
              unloadMuxOut[31] = fifoOut[38][12][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[39][12][w-1];
              unloadMuxOut[1] = fifoOut[40][12][w-1];
              unloadMuxOut[2] = fifoOut[41][12][w-1];
              unloadMuxOut[3] = fifoOut[42][12][w-1];
              unloadMuxOut[4] = fifoOut[43][12][w-1];
              unloadMuxOut[5] = fifoOut[44][12][w-1];
              unloadMuxOut[6] = fifoOut[45][12][w-1];
              unloadMuxOut[7] = fifoOut[46][12][w-1];
              unloadMuxOut[8] = fifoOut[47][12][w-1];
              unloadMuxOut[9] = fifoOut[48][12][w-1];
              unloadMuxOut[10] = fifoOut[49][12][w-1];
              unloadMuxOut[11] = fifoOut[50][12][w-1];
              unloadMuxOut[12] = fifoOut[51][12][w-1];
              unloadMuxOut[13] = fifoOut[26][11][w-1];
              unloadMuxOut[14] = fifoOut[27][11][w-1];
              unloadMuxOut[15] = fifoOut[28][11][w-1];
              unloadMuxOut[16] = fifoOut[29][11][w-1];
              unloadMuxOut[17] = fifoOut[30][11][w-1];
              unloadMuxOut[18] = fifoOut[31][11][w-1];
              unloadMuxOut[19] = fifoOut[32][11][w-1];
              unloadMuxOut[20] = fifoOut[33][11][w-1];
              unloadMuxOut[21] = fifoOut[34][11][w-1];
              unloadMuxOut[22] = fifoOut[35][11][w-1];
              unloadMuxOut[23] = fifoOut[36][11][w-1];
              unloadMuxOut[24] = fifoOut[37][11][w-1];
              unloadMuxOut[25] = fifoOut[38][11][w-1];
              unloadMuxOut[26] = fifoOut[39][11][w-1];
              unloadMuxOut[27] = fifoOut[40][11][w-1];
              unloadMuxOut[28] = fifoOut[41][11][w-1];
              unloadMuxOut[29] = fifoOut[42][11][w-1];
              unloadMuxOut[30] = fifoOut[43][11][w-1];
              unloadMuxOut[31] = fifoOut[44][11][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[45][11][w-1];
              unloadMuxOut[1] = fifoOut[46][11][w-1];
              unloadMuxOut[2] = fifoOut[47][11][w-1];
              unloadMuxOut[3] = fifoOut[48][11][w-1];
              unloadMuxOut[4] = fifoOut[49][11][w-1];
              unloadMuxOut[5] = fifoOut[50][11][w-1];
              unloadMuxOut[6] = fifoOut[51][11][w-1];
              unloadMuxOut[7] = fifoOut[26][10][w-1];
              unloadMuxOut[8] = fifoOut[27][10][w-1];
              unloadMuxOut[9] = fifoOut[28][10][w-1];
              unloadMuxOut[10] = fifoOut[29][10][w-1];
              unloadMuxOut[11] = fifoOut[30][10][w-1];
              unloadMuxOut[12] = fifoOut[31][10][w-1];
              unloadMuxOut[13] = fifoOut[32][10][w-1];
              unloadMuxOut[14] = fifoOut[33][10][w-1];
              unloadMuxOut[15] = fifoOut[34][10][w-1];
              unloadMuxOut[16] = fifoOut[35][10][w-1];
              unloadMuxOut[17] = fifoOut[36][10][w-1];
              unloadMuxOut[18] = fifoOut[37][10][w-1];
              unloadMuxOut[19] = fifoOut[38][10][w-1];
              unloadMuxOut[20] = fifoOut[39][10][w-1];
              unloadMuxOut[21] = fifoOut[40][10][w-1];
              unloadMuxOut[22] = fifoOut[41][10][w-1];
              unloadMuxOut[23] = fifoOut[42][10][w-1];
              unloadMuxOut[24] = fifoOut[43][10][w-1];
              unloadMuxOut[25] = fifoOut[44][10][w-1];
              unloadMuxOut[26] = fifoOut[45][10][w-1];
              unloadMuxOut[27] = fifoOut[46][10][w-1];
              unloadMuxOut[28] = fifoOut[47][10][w-1];
              unloadMuxOut[29] = fifoOut[48][10][w-1];
              unloadMuxOut[30] = fifoOut[49][10][w-1];
              unloadMuxOut[31] = fifoOut[50][10][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[51][10][w-1];
              unloadMuxOut[1] = fifoOut[26][9][w-1];
              unloadMuxOut[2] = fifoOut[27][9][w-1];
              unloadMuxOut[3] = fifoOut[28][9][w-1];
              unloadMuxOut[4] = fifoOut[29][9][w-1];
              unloadMuxOut[5] = fifoOut[30][9][w-1];
              unloadMuxOut[6] = fifoOut[31][9][w-1];
              unloadMuxOut[7] = fifoOut[32][9][w-1];
              unloadMuxOut[8] = fifoOut[33][9][w-1];
              unloadMuxOut[9] = fifoOut[34][9][w-1];
              unloadMuxOut[10] = fifoOut[35][9][w-1];
              unloadMuxOut[11] = fifoOut[36][9][w-1];
              unloadMuxOut[12] = fifoOut[37][9][w-1];
              unloadMuxOut[13] = fifoOut[38][9][w-1];
              unloadMuxOut[14] = fifoOut[39][9][w-1];
              unloadMuxOut[15] = fifoOut[40][9][w-1];
              unloadMuxOut[16] = fifoOut[41][9][w-1];
              unloadMuxOut[17] = fifoOut[42][9][w-1];
              unloadMuxOut[18] = fifoOut[43][9][w-1];
              unloadMuxOut[19] = fifoOut[44][9][w-1];
              unloadMuxOut[20] = fifoOut[45][9][w-1];
              unloadMuxOut[21] = fifoOut[46][9][w-1];
              unloadMuxOut[22] = fifoOut[47][9][w-1];
              unloadMuxOut[23] = fifoOut[48][9][w-1];
              unloadMuxOut[24] = fifoOut[49][9][w-1];
              unloadMuxOut[25] = fifoOut[50][9][w-1];
              unloadMuxOut[26] = fifoOut[51][9][w-1];
              unloadMuxOut[27] = fifoOut[26][8][w-1];
              unloadMuxOut[28] = fifoOut[27][8][w-1];
              unloadMuxOut[29] = fifoOut[28][8][w-1];
              unloadMuxOut[30] = fifoOut[29][8][w-1];
              unloadMuxOut[31] = fifoOut[30][8][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[31][8][w-1];
              unloadMuxOut[1] = fifoOut[32][8][w-1];
              unloadMuxOut[2] = fifoOut[33][8][w-1];
              unloadMuxOut[3] = fifoOut[34][8][w-1];
              unloadMuxOut[4] = fifoOut[35][8][w-1];
              unloadMuxOut[5] = fifoOut[36][8][w-1];
              unloadMuxOut[6] = fifoOut[37][8][w-1];
              unloadMuxOut[7] = fifoOut[38][8][w-1];
              unloadMuxOut[8] = fifoOut[39][8][w-1];
              unloadMuxOut[9] = fifoOut[40][8][w-1];
              unloadMuxOut[10] = fifoOut[41][8][w-1];
              unloadMuxOut[11] = fifoOut[42][8][w-1];
              unloadMuxOut[12] = fifoOut[43][8][w-1];
              unloadMuxOut[13] = fifoOut[44][8][w-1];
              unloadMuxOut[14] = fifoOut[45][8][w-1];
              unloadMuxOut[15] = fifoOut[46][8][w-1];
              unloadMuxOut[16] = fifoOut[47][8][w-1];
              unloadMuxOut[17] = fifoOut[48][8][w-1];
              unloadMuxOut[18] = fifoOut[49][8][w-1];
              unloadMuxOut[19] = fifoOut[50][8][w-1];
              unloadMuxOut[20] = fifoOut[51][8][w-1];
              unloadMuxOut[21] = fifoOut[26][7][w-1];
              unloadMuxOut[22] = fifoOut[27][7][w-1];
              unloadMuxOut[23] = fifoOut[28][7][w-1];
              unloadMuxOut[24] = fifoOut[29][7][w-1];
              unloadMuxOut[25] = fifoOut[30][7][w-1];
              unloadMuxOut[26] = fifoOut[31][7][w-1];
              unloadMuxOut[27] = fifoOut[32][7][w-1];
              unloadMuxOut[28] = fifoOut[33][7][w-1];
              unloadMuxOut[29] = fifoOut[34][7][w-1];
              unloadMuxOut[30] = fifoOut[35][7][w-1];
              unloadMuxOut[31] = fifoOut[36][7][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[37][7][w-1];
              unloadMuxOut[1] = fifoOut[38][7][w-1];
              unloadMuxOut[2] = fifoOut[39][7][w-1];
              unloadMuxOut[3] = fifoOut[40][7][w-1];
              unloadMuxOut[4] = fifoOut[41][7][w-1];
              unloadMuxOut[5] = fifoOut[42][7][w-1];
              unloadMuxOut[6] = fifoOut[43][7][w-1];
              unloadMuxOut[7] = fifoOut[44][7][w-1];
              unloadMuxOut[8] = fifoOut[45][7][w-1];
              unloadMuxOut[9] = fifoOut[46][7][w-1];
              unloadMuxOut[10] = fifoOut[47][7][w-1];
              unloadMuxOut[11] = fifoOut[48][7][w-1];
              unloadMuxOut[12] = fifoOut[49][7][w-1];
              unloadMuxOut[13] = fifoOut[50][7][w-1];
              unloadMuxOut[14] = fifoOut[51][7][w-1];
              unloadMuxOut[15] = fifoOut[26][6][w-1];
              unloadMuxOut[16] = fifoOut[27][6][w-1];
              unloadMuxOut[17] = fifoOut[28][6][w-1];
              unloadMuxOut[18] = fifoOut[29][6][w-1];
              unloadMuxOut[19] = fifoOut[30][6][w-1];
              unloadMuxOut[20] = fifoOut[31][6][w-1];
              unloadMuxOut[21] = fifoOut[32][6][w-1];
              unloadMuxOut[22] = fifoOut[33][6][w-1];
              unloadMuxOut[23] = fifoOut[34][6][w-1];
              unloadMuxOut[24] = fifoOut[35][6][w-1];
              unloadMuxOut[25] = fifoOut[36][6][w-1];
              unloadMuxOut[26] = fifoOut[37][6][w-1];
              unloadMuxOut[27] = fifoOut[38][6][w-1];
              unloadMuxOut[28] = fifoOut[39][6][w-1];
              unloadMuxOut[29] = fifoOut[40][6][w-1];
              unloadMuxOut[30] = fifoOut[41][6][w-1];
              unloadMuxOut[31] = fifoOut[42][6][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[43][6][w-1];
              unloadMuxOut[1] = fifoOut[44][6][w-1];
              unloadMuxOut[2] = fifoOut[45][6][w-1];
              unloadMuxOut[3] = fifoOut[46][6][w-1];
              unloadMuxOut[4] = fifoOut[47][6][w-1];
              unloadMuxOut[5] = fifoOut[48][6][w-1];
              unloadMuxOut[6] = fifoOut[49][6][w-1];
              unloadMuxOut[7] = fifoOut[50][6][w-1];
              unloadMuxOut[8] = fifoOut[51][6][w-1];
              unloadMuxOut[9] = fifoOut[26][5][w-1];
              unloadMuxOut[10] = fifoOut[27][5][w-1];
              unloadMuxOut[11] = fifoOut[28][5][w-1];
              unloadMuxOut[12] = fifoOut[29][5][w-1];
              unloadMuxOut[13] = fifoOut[30][5][w-1];
              unloadMuxOut[14] = fifoOut[31][5][w-1];
              unloadMuxOut[15] = fifoOut[32][5][w-1];
              unloadMuxOut[16] = fifoOut[33][5][w-1];
              unloadMuxOut[17] = fifoOut[34][5][w-1];
              unloadMuxOut[18] = fifoOut[35][5][w-1];
              unloadMuxOut[19] = fifoOut[36][5][w-1];
              unloadMuxOut[20] = fifoOut[37][5][w-1];
              unloadMuxOut[21] = fifoOut[38][5][w-1];
              unloadMuxOut[22] = fifoOut[39][5][w-1];
              unloadMuxOut[23] = fifoOut[40][5][w-1];
              unloadMuxOut[24] = fifoOut[41][5][w-1];
              unloadMuxOut[25] = fifoOut[42][5][w-1];
              unloadMuxOut[26] = fifoOut[43][5][w-1];
              unloadMuxOut[27] = fifoOut[44][5][w-1];
              unloadMuxOut[28] = fifoOut[45][5][w-1];
              unloadMuxOut[29] = fifoOut[46][5][w-1];
              unloadMuxOut[30] = fifoOut[47][5][w-1];
              unloadMuxOut[31] = fifoOut[48][5][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[49][5][w-1];
              unloadMuxOut[1] = fifoOut[50][5][w-1];
              unloadMuxOut[2] = fifoOut[51][5][w-1];
              unloadMuxOut[3] = fifoOut[26][4][w-1];
              unloadMuxOut[4] = fifoOut[27][4][w-1];
              unloadMuxOut[5] = fifoOut[28][4][w-1];
              unloadMuxOut[6] = fifoOut[29][4][w-1];
              unloadMuxOut[7] = fifoOut[30][4][w-1];
              unloadMuxOut[8] = fifoOut[31][4][w-1];
              unloadMuxOut[9] = fifoOut[32][4][w-1];
              unloadMuxOut[10] = fifoOut[33][4][w-1];
              unloadMuxOut[11] = fifoOut[34][4][w-1];
              unloadMuxOut[12] = fifoOut[35][4][w-1];
              unloadMuxOut[13] = fifoOut[36][4][w-1];
              unloadMuxOut[14] = fifoOut[37][4][w-1];
              unloadMuxOut[15] = fifoOut[38][4][w-1];
              unloadMuxOut[16] = fifoOut[39][4][w-1];
              unloadMuxOut[17] = fifoOut[40][4][w-1];
              unloadMuxOut[18] = fifoOut[41][4][w-1];
              unloadMuxOut[19] = fifoOut[42][4][w-1];
              unloadMuxOut[20] = fifoOut[43][4][w-1];
              unloadMuxOut[21] = fifoOut[44][4][w-1];
              unloadMuxOut[22] = fifoOut[45][4][w-1];
              unloadMuxOut[23] = fifoOut[46][4][w-1];
              unloadMuxOut[24] = fifoOut[47][4][w-1];
              unloadMuxOut[25] = fifoOut[48][4][w-1];
              unloadMuxOut[26] = fifoOut[49][4][w-1];
              unloadMuxOut[27] = fifoOut[50][4][w-1];
              unloadMuxOut[28] = fifoOut[51][4][w-1];
              unloadMuxOut[29] = fifoOut[26][3][w-1];
              unloadMuxOut[30] = fifoOut[27][3][w-1];
              unloadMuxOut[31] = fifoOut[28][3][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[29][3][w-1];
              unloadMuxOut[1] = fifoOut[30][3][w-1];
              unloadMuxOut[2] = fifoOut[31][3][w-1];
              unloadMuxOut[3] = fifoOut[32][3][w-1];
              unloadMuxOut[4] = fifoOut[33][3][w-1];
              unloadMuxOut[5] = fifoOut[34][3][w-1];
              unloadMuxOut[6] = fifoOut[35][3][w-1];
              unloadMuxOut[7] = fifoOut[36][3][w-1];
              unloadMuxOut[8] = fifoOut[37][3][w-1];
              unloadMuxOut[9] = fifoOut[38][3][w-1];
              unloadMuxOut[10] = fifoOut[39][3][w-1];
              unloadMuxOut[11] = fifoOut[40][3][w-1];
              unloadMuxOut[12] = fifoOut[41][3][w-1];
              unloadMuxOut[13] = fifoOut[42][3][w-1];
              unloadMuxOut[14] = fifoOut[43][3][w-1];
              unloadMuxOut[15] = fifoOut[44][3][w-1];
              unloadMuxOut[16] = fifoOut[45][3][w-1];
              unloadMuxOut[17] = fifoOut[46][3][w-1];
              unloadMuxOut[18] = fifoOut[47][3][w-1];
              unloadMuxOut[19] = fifoOut[48][3][w-1];
              unloadMuxOut[20] = fifoOut[49][3][w-1];
              unloadMuxOut[21] = fifoOut[50][3][w-1];
              unloadMuxOut[22] = fifoOut[51][3][w-1];
              unloadMuxOut[23] = fifoOut[26][2][w-1];
              unloadMuxOut[24] = fifoOut[27][2][w-1];
              unloadMuxOut[25] = fifoOut[28][2][w-1];
              unloadMuxOut[26] = fifoOut[29][2][w-1];
              unloadMuxOut[27] = fifoOut[30][2][w-1];
              unloadMuxOut[28] = fifoOut[31][2][w-1];
              unloadMuxOut[29] = fifoOut[32][2][w-1];
              unloadMuxOut[30] = fifoOut[33][2][w-1];
              unloadMuxOut[31] = fifoOut[34][2][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[35][2][w-1];
              unloadMuxOut[1] = fifoOut[36][2][w-1];
              unloadMuxOut[2] = fifoOut[37][2][w-1];
              unloadMuxOut[3] = fifoOut[38][2][w-1];
              unloadMuxOut[4] = fifoOut[39][2][w-1];
              unloadMuxOut[5] = fifoOut[40][2][w-1];
              unloadMuxOut[6] = fifoOut[41][2][w-1];
              unloadMuxOut[7] = fifoOut[42][2][w-1];
              unloadMuxOut[8] = fifoOut[43][2][w-1];
              unloadMuxOut[9] = fifoOut[44][2][w-1];
              unloadMuxOut[10] = fifoOut[45][2][w-1];
              unloadMuxOut[11] = fifoOut[46][2][w-1];
              unloadMuxOut[12] = fifoOut[47][2][w-1];
              unloadMuxOut[13] = fifoOut[48][2][w-1];
              unloadMuxOut[14] = fifoOut[49][2][w-1];
              unloadMuxOut[15] = fifoOut[50][2][w-1];
              unloadMuxOut[16] = fifoOut[51][2][w-1];
              unloadMuxOut[17] = fifoOut[26][1][w-1];
              unloadMuxOut[18] = fifoOut[27][1][w-1];
              unloadMuxOut[19] = fifoOut[28][1][w-1];
              unloadMuxOut[20] = fifoOut[29][1][w-1];
              unloadMuxOut[21] = fifoOut[30][1][w-1];
              unloadMuxOut[22] = fifoOut[31][1][w-1];
              unloadMuxOut[23] = fifoOut[32][1][w-1];
              unloadMuxOut[24] = fifoOut[33][1][w-1];
              unloadMuxOut[25] = fifoOut[34][1][w-1];
              unloadMuxOut[26] = fifoOut[35][1][w-1];
              unloadMuxOut[27] = fifoOut[36][1][w-1];
              unloadMuxOut[28] = fifoOut[37][1][w-1];
              unloadMuxOut[29] = fifoOut[38][1][w-1];
              unloadMuxOut[30] = fifoOut[39][1][w-1];
              unloadMuxOut[31] = fifoOut[40][1][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[41][1][w-1];
              unloadMuxOut[1] = fifoOut[42][1][w-1];
              unloadMuxOut[2] = fifoOut[43][1][w-1];
              unloadMuxOut[3] = fifoOut[44][1][w-1];
              unloadMuxOut[4] = fifoOut[45][1][w-1];
              unloadMuxOut[5] = fifoOut[46][1][w-1];
              unloadMuxOut[6] = fifoOut[47][1][w-1];
              unloadMuxOut[7] = fifoOut[48][1][w-1];
              unloadMuxOut[8] = fifoOut[49][1][w-1];
              unloadMuxOut[9] = fifoOut[50][1][w-1];
              unloadMuxOut[10] = fifoOut[51][1][w-1];
              unloadMuxOut[11] = fifoOut[0][12][w-1];
              unloadMuxOut[12] = fifoOut[1][12][w-1];
              unloadMuxOut[13] = fifoOut[2][12][w-1];
              unloadMuxOut[14] = fifoOut[3][12][w-1];
              unloadMuxOut[15] = fifoOut[4][12][w-1];
              unloadMuxOut[16] = fifoOut[5][12][w-1];
              unloadMuxOut[17] = fifoOut[6][12][w-1];
              unloadMuxOut[18] = fifoOut[7][12][w-1];
              unloadMuxOut[19] = fifoOut[8][12][w-1];
              unloadMuxOut[20] = fifoOut[9][12][w-1];
              unloadMuxOut[21] = fifoOut[10][12][w-1];
              unloadMuxOut[22] = fifoOut[11][12][w-1];
              unloadMuxOut[23] = fifoOut[12][12][w-1];
              unloadMuxOut[24] = fifoOut[13][12][w-1];
              unloadMuxOut[25] = fifoOut[14][12][w-1];
              unloadMuxOut[26] = fifoOut[15][12][w-1];
              unloadMuxOut[27] = fifoOut[16][12][w-1];
              unloadMuxOut[28] = fifoOut[17][12][w-1];
              unloadMuxOut[29] = fifoOut[18][12][w-1];
              unloadMuxOut[30] = fifoOut[19][12][w-1];
              unloadMuxOut[31] = fifoOut[20][12][w-1];
       end
       16: begin
              unloadMuxOut[0] = fifoOut[21][12][w-1];
              unloadMuxOut[1] = fifoOut[22][12][w-1];
              unloadMuxOut[2] = fifoOut[23][12][w-1];
              unloadMuxOut[3] = fifoOut[24][12][w-1];
              unloadMuxOut[4] = fifoOut[25][12][w-1];
              unloadMuxOut[5] = fifoOut[0][11][w-1];
              unloadMuxOut[6] = fifoOut[1][11][w-1];
              unloadMuxOut[7] = fifoOut[2][11][w-1];
              unloadMuxOut[8] = fifoOut[3][11][w-1];
              unloadMuxOut[9] = fifoOut[4][11][w-1];
              unloadMuxOut[10] = fifoOut[5][11][w-1];
              unloadMuxOut[11] = fifoOut[6][11][w-1];
              unloadMuxOut[12] = fifoOut[7][11][w-1];
              unloadMuxOut[13] = fifoOut[8][11][w-1];
              unloadMuxOut[14] = fifoOut[9][11][w-1];
              unloadMuxOut[15] = fifoOut[10][11][w-1];
              unloadMuxOut[16] = fifoOut[11][11][w-1];
              unloadMuxOut[17] = fifoOut[12][11][w-1];
              unloadMuxOut[18] = fifoOut[13][11][w-1];
              unloadMuxOut[19] = fifoOut[14][11][w-1];
              unloadMuxOut[20] = fifoOut[15][11][w-1];
              unloadMuxOut[21] = fifoOut[16][11][w-1];
              unloadMuxOut[22] = fifoOut[17][11][w-1];
              unloadMuxOut[23] = fifoOut[18][11][w-1];
              unloadMuxOut[24] = fifoOut[19][11][w-1];
              unloadMuxOut[25] = fifoOut[20][11][w-1];
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0;
             end
       end
    endcase
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[16][5];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[49][3];
              muxOutConnector[27] = fifoOut[50][3];
              muxOutConnector[28] = fifoOut[51][3];
              muxOutConnector[29] = fifoOut[26][2];
              muxOutConnector[30] = fifoOut[27][2];
              muxOutConnector[31] = fifoOut[28][2];
              muxOutConnector[32] = fifoOut[29][2];
              muxOutConnector[33] = fifoOut[30][2];
              muxOutConnector[34] = fifoOut[31][2];
              muxOutConnector[35] = fifoOut[32][2];
              muxOutConnector[36] = fifoOut[33][2];
              muxOutConnector[37] = fifoOut[34][2];
              muxOutConnector[38] = fifoOut[35][2];
              muxOutConnector[39] = fifoOut[36][2];
              muxOutConnector[40] = fifoOut[37][2];
              muxOutConnector[41] = fifoOut[38][2];
              muxOutConnector[42] = fifoOut[39][2];
              muxOutConnector[43] = fifoOut[40][2];
              muxOutConnector[44] = fifoOut[41][2];
              muxOutConnector[45] = fifoOut[42][2];
              muxOutConnector[46] = fifoOut[43][2];
              muxOutConnector[47] = fifoOut[44][2];
              muxOutConnector[48] = fifoOut[45][2];
              muxOutConnector[49] = fifoOut[46][2];
              muxOutConnector[50] = fifoOut[47][2];
              muxOutConnector[51] = fifoOut[48][2];
       end
       1: begin
              muxOutConnector[0] = fifoOut[16][5];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[49][3];
              muxOutConnector[27] = fifoOut[50][3];
              muxOutConnector[28] = fifoOut[51][3];
              muxOutConnector[29] = fifoOut[26][2];
              muxOutConnector[30] = fifoOut[27][2];
              muxOutConnector[31] = fifoOut[28][2];
              muxOutConnector[32] = fifoOut[29][2];
              muxOutConnector[33] = fifoOut[30][2];
              muxOutConnector[34] = fifoOut[31][2];
              muxOutConnector[35] = fifoOut[32][2];
              muxOutConnector[36] = fifoOut[33][2];
              muxOutConnector[37] = fifoOut[34][2];
              muxOutConnector[38] = fifoOut[35][2];
              muxOutConnector[39] = fifoOut[36][2];
              muxOutConnector[40] = fifoOut[37][2];
              muxOutConnector[41] = fifoOut[38][2];
              muxOutConnector[42] = fifoOut[39][2];
              muxOutConnector[43] = fifoOut[40][2];
              muxOutConnector[44] = fifoOut[41][2];
              muxOutConnector[45] = fifoOut[42][2];
              muxOutConnector[46] = fifoOut[43][2];
              muxOutConnector[47] = fifoOut[44][2];
              muxOutConnector[48] = fifoOut[45][2];
              muxOutConnector[49] = fifoOut[46][2];
              muxOutConnector[50] = fifoOut[47][2];
              muxOutConnector[51] = fifoOut[48][2];
       end
       2: begin
              muxOutConnector[0] = fifoOut[16][5];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[49][3];
              muxOutConnector[27] = fifoOut[50][3];
              muxOutConnector[28] = fifoOut[51][3];
              muxOutConnector[29] = fifoOut[26][2];
              muxOutConnector[30] = fifoOut[27][2];
              muxOutConnector[31] = fifoOut[28][2];
              muxOutConnector[32] = fifoOut[29][2];
              muxOutConnector[33] = fifoOut[30][2];
              muxOutConnector[34] = fifoOut[31][2];
              muxOutConnector[35] = fifoOut[32][2];
              muxOutConnector[36] = fifoOut[33][2];
              muxOutConnector[37] = fifoOut[34][2];
              muxOutConnector[38] = fifoOut[35][2];
              muxOutConnector[39] = fifoOut[36][2];
              muxOutConnector[40] = fifoOut[37][2];
              muxOutConnector[41] = fifoOut[38][2];
              muxOutConnector[42] = fifoOut[39][2];
              muxOutConnector[43] = fifoOut[40][2];
              muxOutConnector[44] = fifoOut[41][2];
              muxOutConnector[45] = fifoOut[42][2];
              muxOutConnector[46] = fifoOut[17][1];
              muxOutConnector[47] = fifoOut[18][1];
              muxOutConnector[48] = fifoOut[19][1];
              muxOutConnector[49] = fifoOut[20][1];
              muxOutConnector[50] = fifoOut[21][1];
              muxOutConnector[51] = fifoOut[22][1];
       end
       3: begin
              muxOutConnector[0] = fifoOut[16][5];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[23][2];
              muxOutConnector[27] = fifoOut[24][2];
              muxOutConnector[28] = fifoOut[25][2];
              muxOutConnector[29] = fifoOut[0][1];
              muxOutConnector[30] = fifoOut[1][1];
              muxOutConnector[31] = fifoOut[2][1];
              muxOutConnector[32] = fifoOut[3][1];
              muxOutConnector[33] = fifoOut[4][1];
              muxOutConnector[34] = fifoOut[5][1];
              muxOutConnector[35] = fifoOut[6][1];
              muxOutConnector[36] = fifoOut[7][1];
              muxOutConnector[37] = fifoOut[8][1];
              muxOutConnector[38] = fifoOut[9][1];
              muxOutConnector[39] = fifoOut[10][1];
              muxOutConnector[40] = fifoOut[11][1];
              muxOutConnector[41] = fifoOut[12][1];
              muxOutConnector[42] = fifoOut[13][1];
              muxOutConnector[43] = fifoOut[14][1];
              muxOutConnector[44] = fifoOut[15][1];
              muxOutConnector[45] = fifoOut[16][1];
              muxOutConnector[46] = fifoOut[17][1];
              muxOutConnector[47] = fifoOut[18][1];
              muxOutConnector[48] = fifoOut[19][1];
              muxOutConnector[49] = fifoOut[20][1];
              muxOutConnector[50] = fifoOut[21][1];
              muxOutConnector[51] = fifoOut[22][1];
       end
       4: begin
              muxOutConnector[0] = fifoOut[16][5];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[23][2];
              muxOutConnector[27] = fifoOut[24][2];
              muxOutConnector[28] = fifoOut[25][2];
              muxOutConnector[29] = fifoOut[0][1];
              muxOutConnector[30] = fifoOut[1][1];
              muxOutConnector[31] = fifoOut[2][1];
              muxOutConnector[32] = fifoOut[3][1];
              muxOutConnector[33] = fifoOut[4][1];
              muxOutConnector[34] = fifoOut[5][1];
              muxOutConnector[35] = fifoOut[6][1];
              muxOutConnector[36] = fifoOut[7][1];
              muxOutConnector[37] = fifoOut[8][1];
              muxOutConnector[38] = fifoOut[9][1];
              muxOutConnector[39] = fifoOut[10][1];
              muxOutConnector[40] = fifoOut[11][1];
              muxOutConnector[41] = fifoOut[12][1];
              muxOutConnector[42] = fifoOut[13][1];
              muxOutConnector[43] = fifoOut[14][1];
              muxOutConnector[44] = fifoOut[15][1];
              muxOutConnector[45] = fifoOut[16][1];
              muxOutConnector[46] = fifoOut[17][1];
              muxOutConnector[47] = fifoOut[18][1];
              muxOutConnector[48] = fifoOut[19][1];
              muxOutConnector[49] = fifoOut[20][1];
              muxOutConnector[50] = fifoOut[21][1];
              muxOutConnector[51] = fifoOut[22][1];
       end
       5: begin
              muxOutConnector[0] = fifoOut[16][5];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[23][2];
              muxOutConnector[27] = fifoOut[24][2];
              muxOutConnector[28] = fifoOut[25][2];
              muxOutConnector[29] = fifoOut[0][1];
              muxOutConnector[30] = fifoOut[1][1];
              muxOutConnector[31] = fifoOut[2][1];
              muxOutConnector[32] = fifoOut[3][1];
              muxOutConnector[33] = fifoOut[4][1];
              muxOutConnector[34] = fifoOut[5][1];
              muxOutConnector[35] = fifoOut[6][1];
              muxOutConnector[36] = fifoOut[7][1];
              muxOutConnector[37] = fifoOut[8][1];
              muxOutConnector[38] = fifoOut[9][1];
              muxOutConnector[39] = fifoOut[10][1];
              muxOutConnector[40] = fifoOut[11][1];
              muxOutConnector[41] = fifoOut[12][1];
              muxOutConnector[42] = fifoOut[13][1];
              muxOutConnector[43] = fifoOut[14][1];
              muxOutConnector[44] = fifoOut[15][1];
              muxOutConnector[45] = fifoOut[16][1];
              muxOutConnector[46] = fifoOut[17][1];
              muxOutConnector[47] = fifoOut[18][1];
              muxOutConnector[48] = fifoOut[19][1];
              muxOutConnector[49] = fifoOut[20][1];
              muxOutConnector[50] = fifoOut[21][1];
              muxOutConnector[51] = fifoOut[22][1];
       end
       6: begin
              muxOutConnector[0] = fifoOut[51][0];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[23][2];
              muxOutConnector[27] = fifoOut[24][2];
              muxOutConnector[28] = fifoOut[25][2];
              muxOutConnector[29] = fifoOut[0][1];
              muxOutConnector[30] = fifoOut[1][1];
              muxOutConnector[31] = fifoOut[2][1];
              muxOutConnector[32] = fifoOut[3][1];
              muxOutConnector[33] = fifoOut[4][1];
              muxOutConnector[34] = fifoOut[5][1];
              muxOutConnector[35] = fifoOut[6][1];
              muxOutConnector[36] = fifoOut[7][1];
              muxOutConnector[37] = fifoOut[8][1];
              muxOutConnector[38] = fifoOut[9][1];
              muxOutConnector[39] = fifoOut[10][1];
              muxOutConnector[40] = fifoOut[11][1];
              muxOutConnector[41] = fifoOut[12][1];
              muxOutConnector[42] = fifoOut[13][1];
              muxOutConnector[43] = fifoOut[14][1];
              muxOutConnector[44] = fifoOut[15][1];
              muxOutConnector[45] = fifoOut[16][1];
              muxOutConnector[46] = fifoOut[17][1];
              muxOutConnector[47] = fifoOut[18][1];
              muxOutConnector[48] = fifoOut[19][1];
              muxOutConnector[49] = fifoOut[20][1];
              muxOutConnector[50] = fifoOut[21][1];
              muxOutConnector[51] = fifoOut[22][1];
       end
       7: begin
              muxOutConnector[0] = fifoOut[51][0];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[23][2];
              muxOutConnector[27] = fifoOut[24][2];
              muxOutConnector[28] = fifoOut[25][2];
              muxOutConnector[29] = fifoOut[0][1];
              muxOutConnector[30] = fifoOut[1][1];
              muxOutConnector[31] = fifoOut[2][1];
              muxOutConnector[32] = fifoOut[3][1];
              muxOutConnector[33] = fifoOut[4][1];
              muxOutConnector[34] = fifoOut[5][1];
              muxOutConnector[35] = fifoOut[6][1];
              muxOutConnector[36] = fifoOut[7][1];
              muxOutConnector[37] = fifoOut[8][1];
              muxOutConnector[38] = fifoOut[9][1];
              muxOutConnector[39] = fifoOut[10][1];
              muxOutConnector[40] = fifoOut[11][1];
              muxOutConnector[41] = fifoOut[12][1];
              muxOutConnector[42] = fifoOut[13][1];
              muxOutConnector[43] = fifoOut[14][1];
              muxOutConnector[44] = fifoOut[15][1];
              muxOutConnector[45] = fifoOut[16][1];
              muxOutConnector[46] = fifoOut[17][1];
              muxOutConnector[47] = fifoOut[18][1];
              muxOutConnector[48] = fifoOut[19][1];
              muxOutConnector[49] = fifoOut[20][1];
              muxOutConnector[50] = fifoOut[21][1];
              muxOutConnector[51] = fifoOut[22][1];
       end
       8: begin
              muxOutConnector[0] = fifoOut[51][0];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[23][2];
              muxOutConnector[27] = fifoOut[24][2];
              muxOutConnector[28] = fifoOut[25][2];
              muxOutConnector[29] = fifoOut[0][1];
              muxOutConnector[30] = fifoOut[1][1];
              muxOutConnector[31] = fifoOut[2][1];
              muxOutConnector[32] = fifoOut[3][1];
              muxOutConnector[33] = fifoOut[4][1];
              muxOutConnector[34] = fifoOut[5][1];
              muxOutConnector[35] = fifoOut[6][1];
              muxOutConnector[36] = fifoOut[7][1];
              muxOutConnector[37] = fifoOut[8][1];
              muxOutConnector[38] = fifoOut[9][1];
              muxOutConnector[39] = fifoOut[10][1];
              muxOutConnector[40] = fifoOut[11][1];
              muxOutConnector[41] = fifoOut[12][1];
              muxOutConnector[42] = fifoOut[13][1];
              muxOutConnector[43] = fifoOut[14][1];
              muxOutConnector[44] = fifoOut[15][1];
              muxOutConnector[45] = fifoOut[16][1];
              muxOutConnector[46] = fifoOut[17][1];
              muxOutConnector[47] = fifoOut[18][1];
              muxOutConnector[48] = fifoOut[19][1];
              muxOutConnector[49] = fifoOut[20][1];
              muxOutConnector[50] = fifoOut[21][1];
              muxOutConnector[51] = fifoOut[22][1];
       end
       9: begin
              muxOutConnector[0] = fifoOut[51][0];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[23][2];
              muxOutConnector[27] = fifoOut[24][2];
              muxOutConnector[28] = fifoOut[25][2];
              muxOutConnector[29] = fifoOut[0][1];
              muxOutConnector[30] = fifoOut[1][1];
              muxOutConnector[31] = fifoOut[2][1];
              muxOutConnector[32] = fifoOut[3][1];
              muxOutConnector[33] = fifoOut[4][1];
              muxOutConnector[34] = fifoOut[5][1];
              muxOutConnector[35] = fifoOut[6][1];
              muxOutConnector[36] = fifoOut[7][1];
              muxOutConnector[37] = fifoOut[8][1];
              muxOutConnector[38] = fifoOut[9][1];
              muxOutConnector[39] = fifoOut[10][1];
              muxOutConnector[40] = fifoOut[11][1];
              muxOutConnector[41] = fifoOut[12][1];
              muxOutConnector[42] = fifoOut[13][1];
              muxOutConnector[43] = fifoOut[14][1];
              muxOutConnector[44] = fifoOut[15][1];
              muxOutConnector[45] = fifoOut[16][1];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       10: begin
              muxOutConnector[0] = fifoOut[51][0];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       11: begin
              muxOutConnector[0] = fifoOut[51][0];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       12: begin
              muxOutConnector[0] = fifoOut[51][0];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[17][11];
              muxOutConnector[19] = fifoOut[18][11];
              muxOutConnector[20] = fifoOut[19][11];
              muxOutConnector[21] = fifoOut[20][11];
              muxOutConnector[22] = fifoOut[21][11];
              muxOutConnector[23] = fifoOut[22][11];
              muxOutConnector[24] = fifoOut[23][11];
              muxOutConnector[25] = fifoOut[24][11];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       13: begin
              muxOutConnector[0] = fifoOut[25][12];
              muxOutConnector[1] = fifoOut[0][11];
              muxOutConnector[2] = fifoOut[1][11];
              muxOutConnector[3] = fifoOut[2][11];
              muxOutConnector[4] = fifoOut[3][11];
              muxOutConnector[5] = fifoOut[4][11];
              muxOutConnector[6] = fifoOut[5][11];
              muxOutConnector[7] = fifoOut[6][11];
              muxOutConnector[8] = fifoOut[7][11];
              muxOutConnector[9] = fifoOut[8][11];
              muxOutConnector[10] = fifoOut[9][11];
              muxOutConnector[11] = fifoOut[10][11];
              muxOutConnector[12] = fifoOut[11][11];
              muxOutConnector[13] = fifoOut[12][11];
              muxOutConnector[14] = fifoOut[13][11];
              muxOutConnector[15] = fifoOut[14][11];
              muxOutConnector[16] = fifoOut[15][11];
              muxOutConnector[17] = fifoOut[16][11];
              muxOutConnector[18] = fifoOut[17][11];
              muxOutConnector[19] = fifoOut[18][11];
              muxOutConnector[20] = fifoOut[19][11];
              muxOutConnector[21] = fifoOut[20][11];
              muxOutConnector[22] = fifoOut[21][11];
              muxOutConnector[23] = fifoOut[22][11];
              muxOutConnector[24] = fifoOut[23][11];
              muxOutConnector[25] = fifoOut[24][11];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       14: begin
              muxOutConnector[0] = fifoOut[25][12];
              muxOutConnector[1] = fifoOut[0][11];
              muxOutConnector[2] = fifoOut[1][11];
              muxOutConnector[3] = fifoOut[2][11];
              muxOutConnector[4] = fifoOut[3][11];
              muxOutConnector[5] = fifoOut[4][11];
              muxOutConnector[6] = fifoOut[5][11];
              muxOutConnector[7] = fifoOut[6][11];
              muxOutConnector[8] = fifoOut[7][11];
              muxOutConnector[9] = fifoOut[8][11];
              muxOutConnector[10] = fifoOut[9][11];
              muxOutConnector[11] = fifoOut[10][11];
              muxOutConnector[12] = fifoOut[11][11];
              muxOutConnector[13] = fifoOut[12][11];
              muxOutConnector[14] = fifoOut[13][11];
              muxOutConnector[15] = fifoOut[14][11];
              muxOutConnector[16] = fifoOut[15][11];
              muxOutConnector[17] = fifoOut[16][11];
              muxOutConnector[18] = fifoOut[17][11];
              muxOutConnector[19] = fifoOut[18][11];
              muxOutConnector[20] = fifoOut[19][11];
              muxOutConnector[21] = fifoOut[20][11];
              muxOutConnector[22] = fifoOut[21][11];
              muxOutConnector[23] = fifoOut[22][11];
              muxOutConnector[24] = fifoOut[23][11];
              muxOutConnector[25] = fifoOut[24][11];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       15: begin
              muxOutConnector[0] = fifoOut[25][12];
              muxOutConnector[1] = fifoOut[0][11];
              muxOutConnector[2] = fifoOut[1][11];
              muxOutConnector[3] = fifoOut[2][11];
              muxOutConnector[4] = fifoOut[3][11];
              muxOutConnector[5] = fifoOut[4][11];
              muxOutConnector[6] = fifoOut[5][11];
              muxOutConnector[7] = fifoOut[6][11];
              muxOutConnector[8] = fifoOut[7][11];
              muxOutConnector[9] = fifoOut[8][11];
              muxOutConnector[10] = fifoOut[9][11];
              muxOutConnector[11] = fifoOut[10][11];
              muxOutConnector[12] = fifoOut[11][11];
              muxOutConnector[13] = fifoOut[12][11];
              muxOutConnector[14] = fifoOut[13][11];
              muxOutConnector[15] = fifoOut[14][11];
              muxOutConnector[16] = fifoOut[15][11];
              muxOutConnector[17] = fifoOut[16][11];
              muxOutConnector[18] = fifoOut[17][11];
              muxOutConnector[19] = fifoOut[18][11];
              muxOutConnector[20] = fifoOut[19][11];
              muxOutConnector[21] = fifoOut[20][11];
              muxOutConnector[22] = fifoOut[21][11];
              muxOutConnector[23] = fifoOut[22][11];
              muxOutConnector[24] = fifoOut[23][11];
              muxOutConnector[25] = fifoOut[24][11];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       16: begin
              muxOutConnector[0] = fifoOut[25][12];
              muxOutConnector[1] = fifoOut[0][11];
              muxOutConnector[2] = fifoOut[1][11];
              muxOutConnector[3] = fifoOut[2][11];
              muxOutConnector[4] = fifoOut[3][11];
              muxOutConnector[5] = fifoOut[4][11];
              muxOutConnector[6] = fifoOut[5][11];
              muxOutConnector[7] = fifoOut[6][11];
              muxOutConnector[8] = fifoOut[7][11];
              muxOutConnector[9] = fifoOut[8][11];
              muxOutConnector[10] = fifoOut[9][11];
              muxOutConnector[11] = fifoOut[10][11];
              muxOutConnector[12] = fifoOut[11][11];
              muxOutConnector[13] = fifoOut[12][11];
              muxOutConnector[14] = fifoOut[13][11];
              muxOutConnector[15] = fifoOut[14][11];
              muxOutConnector[16] = fifoOut[15][11];
              muxOutConnector[17] = fifoOut[16][11];
              muxOutConnector[18] = fifoOut[17][11];
              muxOutConnector[19] = fifoOut[18][11];
              muxOutConnector[20] = fifoOut[19][11];
              muxOutConnector[21] = fifoOut[20][11];
              muxOutConnector[22] = fifoOut[21][11];
              muxOutConnector[23] = fifoOut[22][11];
              muxOutConnector[24] = fifoOut[23][11];
              muxOutConnector[25] = fifoOut[24][11];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       17: begin
              muxOutConnector[0] = fifoOut[25][12];
              muxOutConnector[1] = fifoOut[0][11];
              muxOutConnector[2] = fifoOut[1][11];
              muxOutConnector[3] = fifoOut[2][11];
              muxOutConnector[4] = fifoOut[3][11];
              muxOutConnector[5] = fifoOut[4][11];
              muxOutConnector[6] = fifoOut[5][11];
              muxOutConnector[7] = fifoOut[6][11];
              muxOutConnector[8] = fifoOut[7][11];
              muxOutConnector[9] = fifoOut[8][11];
              muxOutConnector[10] = fifoOut[9][11];
              muxOutConnector[11] = fifoOut[10][11];
              muxOutConnector[12] = fifoOut[11][11];
              muxOutConnector[13] = fifoOut[12][11];
              muxOutConnector[14] = fifoOut[13][11];
              muxOutConnector[15] = fifoOut[14][11];
              muxOutConnector[16] = fifoOut[15][11];
              muxOutConnector[17] = fifoOut[16][11];
              muxOutConnector[18] = fifoOut[17][11];
              muxOutConnector[19] = fifoOut[18][11];
              muxOutConnector[20] = fifoOut[19][11];
              muxOutConnector[21] = fifoOut[20][11];
              muxOutConnector[22] = fifoOut[21][11];
              muxOutConnector[23] = fifoOut[22][11];
              muxOutConnector[24] = fifoOut[23][11];
              muxOutConnector[25] = fifoOut[24][11];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       18: begin
              muxOutConnector[0] = fifoOut[25][12];
              muxOutConnector[1] = fifoOut[0][11];
              muxOutConnector[2] = fifoOut[1][11];
              muxOutConnector[3] = fifoOut[2][11];
              muxOutConnector[4] = fifoOut[3][11];
              muxOutConnector[5] = fifoOut[4][11];
              muxOutConnector[6] = fifoOut[5][11];
              muxOutConnector[7] = fifoOut[6][11];
              muxOutConnector[8] = fifoOut[7][11];
              muxOutConnector[9] = fifoOut[8][11];
              muxOutConnector[10] = fifoOut[9][11];
              muxOutConnector[11] = fifoOut[10][11];
              muxOutConnector[12] = fifoOut[11][11];
              muxOutConnector[13] = fifoOut[12][11];
              muxOutConnector[14] = fifoOut[13][11];
              muxOutConnector[15] = fifoOut[14][11];
              muxOutConnector[16] = fifoOut[15][11];
              muxOutConnector[17] = fifoOut[16][11];
              muxOutConnector[18] = fifoOut[17][11];
              muxOutConnector[19] = fifoOut[18][11];
              muxOutConnector[20] = fifoOut[19][11];
              muxOutConnector[21] = fifoOut[20][11];
              muxOutConnector[22] = fifoOut[21][11];
              muxOutConnector[23] = fifoOut[22][11];
              muxOutConnector[24] = fifoOut[23][11];
              muxOutConnector[25] = fifoOut[24][11];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       19: begin
              muxOutConnector[0] = fifoOut[25][12];
              muxOutConnector[1] = fifoOut[0][11];
              muxOutConnector[2] = fifoOut[1][11];
              muxOutConnector[3] = fifoOut[2][11];
              muxOutConnector[4] = fifoOut[3][11];
              muxOutConnector[5] = fifoOut[4][11];
              muxOutConnector[6] = fifoOut[5][11];
              muxOutConnector[7] = fifoOut[6][11];
              muxOutConnector[8] = fifoOut[7][11];
              muxOutConnector[9] = fifoOut[8][11];
              muxOutConnector[10] = fifoOut[9][11];
              muxOutConnector[11] = fifoOut[10][11];
              muxOutConnector[12] = fifoOut[11][11];
              muxOutConnector[13] = fifoOut[12][11];
              muxOutConnector[14] = fifoOut[13][11];
              muxOutConnector[15] = fifoOut[14][11];
              muxOutConnector[16] = fifoOut[15][11];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
