`timescale 1ns / 1ps
module LMem1To0_511_ns_yu_circ3_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 12;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input [ADDRESSWIDTH-1:0]unloadAddress;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            fifoOut[i][0] <= ly0InConnector[i];
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
       0: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = fifoOut[17][10][w-1];
              unloadMuxOut[12] = fifoOut[18][10][w-1];
              unloadMuxOut[13] = fifoOut[19][10][w-1];
              unloadMuxOut[14] = fifoOut[20][10][w-1];
              unloadMuxOut[15] = fifoOut[21][10][w-1];
              unloadMuxOut[16] = fifoOut[22][10][w-1];
              unloadMuxOut[17] = fifoOut[23][10][w-1];
              unloadMuxOut[18] = fifoOut[24][10][w-1];
              unloadMuxOut[19] = fifoOut[25][10][w-1];
              unloadMuxOut[20] = fifoOut[0][9][w-1];
              unloadMuxOut[21] = fifoOut[1][9][w-1];
              unloadMuxOut[22] = fifoOut[2][9][w-1];
              unloadMuxOut[23] = fifoOut[3][9][w-1];
              unloadMuxOut[24] = fifoOut[4][9][w-1];
              unloadMuxOut[25] = fifoOut[5][9][w-1];
              unloadMuxOut[26] = fifoOut[6][9][w-1];
              unloadMuxOut[27] = fifoOut[7][9][w-1];
              unloadMuxOut[28] = fifoOut[8][9][w-1];
              unloadMuxOut[29] = fifoOut[9][9][w-1];
              unloadMuxOut[30] = fifoOut[10][9][w-1];
              unloadMuxOut[31] = fifoOut[11][9][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[12][9][w-1];
              unloadMuxOut[1] = fifoOut[13][9][w-1];
              unloadMuxOut[2] = fifoOut[14][9][w-1];
              unloadMuxOut[3] = fifoOut[15][9][w-1];
              unloadMuxOut[4] = fifoOut[16][9][w-1];
              unloadMuxOut[5] = fifoOut[17][9][w-1];
              unloadMuxOut[6] = fifoOut[18][9][w-1];
              unloadMuxOut[7] = fifoOut[19][9][w-1];
              unloadMuxOut[8] = fifoOut[20][9][w-1];
              unloadMuxOut[9] = fifoOut[21][9][w-1];
              unloadMuxOut[10] = fifoOut[22][9][w-1];
              unloadMuxOut[11] = fifoOut[23][9][w-1];
              unloadMuxOut[12] = fifoOut[24][9][w-1];
              unloadMuxOut[13] = fifoOut[25][9][w-1];
              unloadMuxOut[14] = fifoOut[0][8][w-1];
              unloadMuxOut[15] = fifoOut[1][8][w-1];
              unloadMuxOut[16] = fifoOut[2][8][w-1];
              unloadMuxOut[17] = fifoOut[3][8][w-1];
              unloadMuxOut[18] = fifoOut[4][8][w-1];
              unloadMuxOut[19] = fifoOut[5][8][w-1];
              unloadMuxOut[20] = fifoOut[6][8][w-1];
              unloadMuxOut[21] = fifoOut[7][8][w-1];
              unloadMuxOut[22] = fifoOut[8][8][w-1];
              unloadMuxOut[23] = fifoOut[9][8][w-1];
              unloadMuxOut[24] = fifoOut[10][8][w-1];
              unloadMuxOut[25] = fifoOut[11][8][w-1];
              unloadMuxOut[26] = fifoOut[12][8][w-1];
              unloadMuxOut[27] = fifoOut[13][8][w-1];
              unloadMuxOut[28] = fifoOut[14][8][w-1];
              unloadMuxOut[29] = fifoOut[15][8][w-1];
              unloadMuxOut[30] = fifoOut[16][8][w-1];
              unloadMuxOut[31] = fifoOut[17][8][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[18][8][w-1];
              unloadMuxOut[1] = fifoOut[19][8][w-1];
              unloadMuxOut[2] = fifoOut[20][8][w-1];
              unloadMuxOut[3] = fifoOut[21][8][w-1];
              unloadMuxOut[4] = fifoOut[22][8][w-1];
              unloadMuxOut[5] = fifoOut[23][8][w-1];
              unloadMuxOut[6] = fifoOut[24][8][w-1];
              unloadMuxOut[7] = fifoOut[25][8][w-1];
              unloadMuxOut[8] = fifoOut[0][7][w-1];
              unloadMuxOut[9] = fifoOut[1][7][w-1];
              unloadMuxOut[10] = fifoOut[2][7][w-1];
              unloadMuxOut[11] = fifoOut[3][7][w-1];
              unloadMuxOut[12] = fifoOut[4][7][w-1];
              unloadMuxOut[13] = fifoOut[5][7][w-1];
              unloadMuxOut[14] = fifoOut[6][7][w-1];
              unloadMuxOut[15] = fifoOut[7][7][w-1];
              unloadMuxOut[16] = fifoOut[8][7][w-1];
              unloadMuxOut[17] = fifoOut[9][7][w-1];
              unloadMuxOut[18] = fifoOut[10][7][w-1];
              unloadMuxOut[19] = fifoOut[11][7][w-1];
              unloadMuxOut[20] = fifoOut[12][7][w-1];
              unloadMuxOut[21] = fifoOut[13][7][w-1];
              unloadMuxOut[22] = fifoOut[14][7][w-1];
              unloadMuxOut[23] = fifoOut[15][7][w-1];
              unloadMuxOut[24] = fifoOut[16][7][w-1];
              unloadMuxOut[25] = fifoOut[17][7][w-1];
              unloadMuxOut[26] = fifoOut[18][7][w-1];
              unloadMuxOut[27] = fifoOut[19][7][w-1];
              unloadMuxOut[28] = fifoOut[20][7][w-1];
              unloadMuxOut[29] = fifoOut[21][7][w-1];
              unloadMuxOut[30] = fifoOut[22][7][w-1];
              unloadMuxOut[31] = fifoOut[23][7][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[24][7][w-1];
              unloadMuxOut[1] = fifoOut[25][7][w-1];
              unloadMuxOut[2] = fifoOut[0][6][w-1];
              unloadMuxOut[3] = fifoOut[1][6][w-1];
              unloadMuxOut[4] = fifoOut[2][6][w-1];
              unloadMuxOut[5] = fifoOut[3][6][w-1];
              unloadMuxOut[6] = fifoOut[4][6][w-1];
              unloadMuxOut[7] = fifoOut[5][6][w-1];
              unloadMuxOut[8] = fifoOut[6][6][w-1];
              unloadMuxOut[9] = fifoOut[7][6][w-1];
              unloadMuxOut[10] = fifoOut[8][6][w-1];
              unloadMuxOut[11] = fifoOut[9][6][w-1];
              unloadMuxOut[12] = fifoOut[10][6][w-1];
              unloadMuxOut[13] = fifoOut[11][6][w-1];
              unloadMuxOut[14] = fifoOut[12][6][w-1];
              unloadMuxOut[15] = fifoOut[13][6][w-1];
              unloadMuxOut[16] = fifoOut[14][6][w-1];
              unloadMuxOut[17] = fifoOut[15][6][w-1];
              unloadMuxOut[18] = fifoOut[16][6][w-1];
              unloadMuxOut[19] = fifoOut[17][6][w-1];
              unloadMuxOut[20] = fifoOut[18][6][w-1];
              unloadMuxOut[21] = fifoOut[19][6][w-1];
              unloadMuxOut[22] = fifoOut[20][6][w-1];
              unloadMuxOut[23] = fifoOut[21][6][w-1];
              unloadMuxOut[24] = fifoOut[22][6][w-1];
              unloadMuxOut[25] = fifoOut[23][6][w-1];
              unloadMuxOut[26] = fifoOut[24][6][w-1];
              unloadMuxOut[27] = fifoOut[25][6][w-1];
              unloadMuxOut[28] = fifoOut[0][5][w-1];
              unloadMuxOut[29] = fifoOut[1][5][w-1];
              unloadMuxOut[30] = fifoOut[2][5][w-1];
              unloadMuxOut[31] = fifoOut[3][5][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[4][5][w-1];
              unloadMuxOut[1] = fifoOut[5][5][w-1];
              unloadMuxOut[2] = fifoOut[6][5][w-1];
              unloadMuxOut[3] = fifoOut[7][5][w-1];
              unloadMuxOut[4] = fifoOut[8][5][w-1];
              unloadMuxOut[5] = fifoOut[9][5][w-1];
              unloadMuxOut[6] = fifoOut[10][5][w-1];
              unloadMuxOut[7] = fifoOut[11][5][w-1];
              unloadMuxOut[8] = fifoOut[12][5][w-1];
              unloadMuxOut[9] = fifoOut[13][5][w-1];
              unloadMuxOut[10] = fifoOut[14][5][w-1];
              unloadMuxOut[11] = fifoOut[15][5][w-1];
              unloadMuxOut[12] = fifoOut[16][5][w-1];
              unloadMuxOut[13] = fifoOut[17][5][w-1];
              unloadMuxOut[14] = fifoOut[18][5][w-1];
              unloadMuxOut[15] = fifoOut[19][5][w-1];
              unloadMuxOut[16] = fifoOut[20][5][w-1];
              unloadMuxOut[17] = fifoOut[21][5][w-1];
              unloadMuxOut[18] = fifoOut[22][5][w-1];
              unloadMuxOut[19] = fifoOut[23][5][w-1];
              unloadMuxOut[20] = fifoOut[24][5][w-1];
              unloadMuxOut[21] = fifoOut[25][5][w-1];
              unloadMuxOut[22] = fifoOut[0][4][w-1];
              unloadMuxOut[23] = fifoOut[1][4][w-1];
              unloadMuxOut[24] = fifoOut[2][4][w-1];
              unloadMuxOut[25] = fifoOut[3][4][w-1];
              unloadMuxOut[26] = fifoOut[4][4][w-1];
              unloadMuxOut[27] = fifoOut[5][4][w-1];
              unloadMuxOut[28] = fifoOut[6][4][w-1];
              unloadMuxOut[29] = fifoOut[7][4][w-1];
              unloadMuxOut[30] = fifoOut[8][4][w-1];
              unloadMuxOut[31] = fifoOut[9][4][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[10][4][w-1];
              unloadMuxOut[1] = fifoOut[11][4][w-1];
              unloadMuxOut[2] = fifoOut[12][4][w-1];
              unloadMuxOut[3] = fifoOut[13][4][w-1];
              unloadMuxOut[4] = fifoOut[14][4][w-1];
              unloadMuxOut[5] = fifoOut[15][4][w-1];
              unloadMuxOut[6] = fifoOut[16][4][w-1];
              unloadMuxOut[7] = fifoOut[17][4][w-1];
              unloadMuxOut[8] = fifoOut[18][4][w-1];
              unloadMuxOut[9] = fifoOut[19][4][w-1];
              unloadMuxOut[10] = fifoOut[20][4][w-1];
              unloadMuxOut[11] = fifoOut[21][4][w-1];
              unloadMuxOut[12] = fifoOut[22][4][w-1];
              unloadMuxOut[13] = fifoOut[23][4][w-1];
              unloadMuxOut[14] = fifoOut[24][4][w-1];
              unloadMuxOut[15] = fifoOut[25][4][w-1];
              unloadMuxOut[16] = fifoOut[0][3][w-1];
              unloadMuxOut[17] = fifoOut[1][3][w-1];
              unloadMuxOut[18] = fifoOut[2][3][w-1];
              unloadMuxOut[19] = fifoOut[3][3][w-1];
              unloadMuxOut[20] = fifoOut[4][3][w-1];
              unloadMuxOut[21] = fifoOut[5][3][w-1];
              unloadMuxOut[22] = fifoOut[6][3][w-1];
              unloadMuxOut[23] = fifoOut[7][3][w-1];
              unloadMuxOut[24] = fifoOut[8][3][w-1];
              unloadMuxOut[25] = fifoOut[9][3][w-1];
              unloadMuxOut[26] = fifoOut[26][11][w-1];
              unloadMuxOut[27] = fifoOut[27][11][w-1];
              unloadMuxOut[28] = fifoOut[28][11][w-1];
              unloadMuxOut[29] = fifoOut[29][11][w-1];
              unloadMuxOut[30] = fifoOut[30][11][w-1];
              unloadMuxOut[31] = fifoOut[31][11][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[32][11][w-1];
              unloadMuxOut[1] = fifoOut[33][11][w-1];
              unloadMuxOut[2] = fifoOut[34][11][w-1];
              unloadMuxOut[3] = fifoOut[35][11][w-1];
              unloadMuxOut[4] = fifoOut[36][11][w-1];
              unloadMuxOut[5] = fifoOut[37][11][w-1];
              unloadMuxOut[6] = fifoOut[38][11][w-1];
              unloadMuxOut[7] = fifoOut[39][11][w-1];
              unloadMuxOut[8] = fifoOut[40][11][w-1];
              unloadMuxOut[9] = fifoOut[41][11][w-1];
              unloadMuxOut[10] = fifoOut[42][11][w-1];
              unloadMuxOut[11] = fifoOut[43][11][w-1];
              unloadMuxOut[12] = fifoOut[44][11][w-1];
              unloadMuxOut[13] = fifoOut[45][11][w-1];
              unloadMuxOut[14] = fifoOut[46][11][w-1];
              unloadMuxOut[15] = fifoOut[47][11][w-1];
              unloadMuxOut[16] = fifoOut[48][11][w-1];
              unloadMuxOut[17] = fifoOut[49][11][w-1];
              unloadMuxOut[18] = fifoOut[50][11][w-1];
              unloadMuxOut[19] = fifoOut[51][11][w-1];
              unloadMuxOut[20] = fifoOut[26][10][w-1];
              unloadMuxOut[21] = fifoOut[27][10][w-1];
              unloadMuxOut[22] = fifoOut[28][10][w-1];
              unloadMuxOut[23] = fifoOut[29][10][w-1];
              unloadMuxOut[24] = fifoOut[30][10][w-1];
              unloadMuxOut[25] = fifoOut[31][10][w-1];
              unloadMuxOut[26] = fifoOut[32][10][w-1];
              unloadMuxOut[27] = fifoOut[33][10][w-1];
              unloadMuxOut[28] = fifoOut[34][10][w-1];
              unloadMuxOut[29] = fifoOut[35][10][w-1];
              unloadMuxOut[30] = fifoOut[36][10][w-1];
              unloadMuxOut[31] = fifoOut[37][10][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[38][10][w-1];
              unloadMuxOut[1] = fifoOut[39][10][w-1];
              unloadMuxOut[2] = fifoOut[40][10][w-1];
              unloadMuxOut[3] = fifoOut[41][10][w-1];
              unloadMuxOut[4] = fifoOut[42][10][w-1];
              unloadMuxOut[5] = fifoOut[43][10][w-1];
              unloadMuxOut[6] = fifoOut[44][10][w-1];
              unloadMuxOut[7] = fifoOut[45][10][w-1];
              unloadMuxOut[8] = fifoOut[46][10][w-1];
              unloadMuxOut[9] = fifoOut[47][10][w-1];
              unloadMuxOut[10] = fifoOut[48][10][w-1];
              unloadMuxOut[11] = fifoOut[49][10][w-1];
              unloadMuxOut[12] = fifoOut[50][10][w-1];
              unloadMuxOut[13] = fifoOut[51][10][w-1];
              unloadMuxOut[14] = fifoOut[26][9][w-1];
              unloadMuxOut[15] = fifoOut[27][9][w-1];
              unloadMuxOut[16] = fifoOut[28][9][w-1];
              unloadMuxOut[17] = fifoOut[29][9][w-1];
              unloadMuxOut[18] = fifoOut[30][9][w-1];
              unloadMuxOut[19] = fifoOut[31][9][w-1];
              unloadMuxOut[20] = fifoOut[32][9][w-1];
              unloadMuxOut[21] = fifoOut[33][9][w-1];
              unloadMuxOut[22] = fifoOut[34][9][w-1];
              unloadMuxOut[23] = fifoOut[35][9][w-1];
              unloadMuxOut[24] = fifoOut[36][9][w-1];
              unloadMuxOut[25] = fifoOut[37][9][w-1];
              unloadMuxOut[26] = fifoOut[38][9][w-1];
              unloadMuxOut[27] = fifoOut[39][9][w-1];
              unloadMuxOut[28] = fifoOut[40][9][w-1];
              unloadMuxOut[29] = fifoOut[41][9][w-1];
              unloadMuxOut[30] = fifoOut[42][9][w-1];
              unloadMuxOut[31] = fifoOut[43][9][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[44][9][w-1];
              unloadMuxOut[1] = fifoOut[45][9][w-1];
              unloadMuxOut[2] = fifoOut[46][9][w-1];
              unloadMuxOut[3] = fifoOut[47][9][w-1];
              unloadMuxOut[4] = fifoOut[48][9][w-1];
              unloadMuxOut[5] = fifoOut[49][9][w-1];
              unloadMuxOut[6] = fifoOut[50][9][w-1];
              unloadMuxOut[7] = fifoOut[51][9][w-1];
              unloadMuxOut[8] = fifoOut[26][8][w-1];
              unloadMuxOut[9] = fifoOut[27][8][w-1];
              unloadMuxOut[10] = fifoOut[28][8][w-1];
              unloadMuxOut[11] = fifoOut[29][8][w-1];
              unloadMuxOut[12] = fifoOut[30][8][w-1];
              unloadMuxOut[13] = fifoOut[31][8][w-1];
              unloadMuxOut[14] = fifoOut[32][8][w-1];
              unloadMuxOut[15] = fifoOut[33][8][w-1];
              unloadMuxOut[16] = fifoOut[34][8][w-1];
              unloadMuxOut[17] = fifoOut[35][8][w-1];
              unloadMuxOut[18] = fifoOut[36][8][w-1];
              unloadMuxOut[19] = fifoOut[37][8][w-1];
              unloadMuxOut[20] = fifoOut[38][8][w-1];
              unloadMuxOut[21] = fifoOut[39][8][w-1];
              unloadMuxOut[22] = fifoOut[40][8][w-1];
              unloadMuxOut[23] = fifoOut[41][8][w-1];
              unloadMuxOut[24] = fifoOut[42][8][w-1];
              unloadMuxOut[25] = fifoOut[43][8][w-1];
              unloadMuxOut[26] = fifoOut[44][8][w-1];
              unloadMuxOut[27] = fifoOut[45][8][w-1];
              unloadMuxOut[28] = fifoOut[46][8][w-1];
              unloadMuxOut[29] = fifoOut[47][8][w-1];
              unloadMuxOut[30] = fifoOut[48][8][w-1];
              unloadMuxOut[31] = fifoOut[49][8][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[50][8][w-1];
              unloadMuxOut[1] = fifoOut[51][8][w-1];
              unloadMuxOut[2] = fifoOut[26][7][w-1];
              unloadMuxOut[3] = fifoOut[27][7][w-1];
              unloadMuxOut[4] = fifoOut[28][7][w-1];
              unloadMuxOut[5] = fifoOut[29][7][w-1];
              unloadMuxOut[6] = fifoOut[30][7][w-1];
              unloadMuxOut[7] = fifoOut[31][7][w-1];
              unloadMuxOut[8] = fifoOut[32][7][w-1];
              unloadMuxOut[9] = fifoOut[33][7][w-1];
              unloadMuxOut[10] = fifoOut[34][7][w-1];
              unloadMuxOut[11] = fifoOut[35][7][w-1];
              unloadMuxOut[12] = fifoOut[36][7][w-1];
              unloadMuxOut[13] = fifoOut[37][7][w-1];
              unloadMuxOut[14] = fifoOut[38][7][w-1];
              unloadMuxOut[15] = fifoOut[39][7][w-1];
              unloadMuxOut[16] = fifoOut[40][7][w-1];
              unloadMuxOut[17] = fifoOut[41][7][w-1];
              unloadMuxOut[18] = fifoOut[42][7][w-1];
              unloadMuxOut[19] = fifoOut[43][7][w-1];
              unloadMuxOut[20] = fifoOut[44][7][w-1];
              unloadMuxOut[21] = fifoOut[45][7][w-1];
              unloadMuxOut[22] = fifoOut[46][7][w-1];
              unloadMuxOut[23] = fifoOut[47][7][w-1];
              unloadMuxOut[24] = fifoOut[48][7][w-1];
              unloadMuxOut[25] = fifoOut[49][7][w-1];
              unloadMuxOut[26] = fifoOut[50][7][w-1];
              unloadMuxOut[27] = fifoOut[51][7][w-1];
              unloadMuxOut[28] = fifoOut[26][6][w-1];
              unloadMuxOut[29] = fifoOut[27][6][w-1];
              unloadMuxOut[30] = fifoOut[28][6][w-1];
              unloadMuxOut[31] = fifoOut[29][6][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[30][6][w-1];
              unloadMuxOut[1] = fifoOut[31][6][w-1];
              unloadMuxOut[2] = fifoOut[32][6][w-1];
              unloadMuxOut[3] = fifoOut[33][6][w-1];
              unloadMuxOut[4] = fifoOut[34][6][w-1];
              unloadMuxOut[5] = fifoOut[35][6][w-1];
              unloadMuxOut[6] = fifoOut[36][6][w-1];
              unloadMuxOut[7] = fifoOut[37][6][w-1];
              unloadMuxOut[8] = fifoOut[38][6][w-1];
              unloadMuxOut[9] = fifoOut[39][6][w-1];
              unloadMuxOut[10] = fifoOut[40][6][w-1];
              unloadMuxOut[11] = fifoOut[41][6][w-1];
              unloadMuxOut[12] = fifoOut[42][6][w-1];
              unloadMuxOut[13] = fifoOut[43][6][w-1];
              unloadMuxOut[14] = fifoOut[44][6][w-1];
              unloadMuxOut[15] = fifoOut[45][6][w-1];
              unloadMuxOut[16] = fifoOut[46][6][w-1];
              unloadMuxOut[17] = fifoOut[47][6][w-1];
              unloadMuxOut[18] = fifoOut[48][6][w-1];
              unloadMuxOut[19] = fifoOut[49][6][w-1];
              unloadMuxOut[20] = fifoOut[50][6][w-1];
              unloadMuxOut[21] = fifoOut[51][6][w-1];
              unloadMuxOut[22] = fifoOut[26][5][w-1];
              unloadMuxOut[23] = fifoOut[27][5][w-1];
              unloadMuxOut[24] = fifoOut[28][5][w-1];
              unloadMuxOut[25] = fifoOut[29][5][w-1];
              unloadMuxOut[26] = fifoOut[30][5][w-1];
              unloadMuxOut[27] = fifoOut[31][5][w-1];
              unloadMuxOut[28] = fifoOut[32][5][w-1];
              unloadMuxOut[29] = fifoOut[33][5][w-1];
              unloadMuxOut[30] = fifoOut[34][5][w-1];
              unloadMuxOut[31] = fifoOut[35][5][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[36][5][w-1];
              unloadMuxOut[1] = fifoOut[37][5][w-1];
              unloadMuxOut[2] = fifoOut[38][5][w-1];
              unloadMuxOut[3] = fifoOut[39][5][w-1];
              unloadMuxOut[4] = fifoOut[40][5][w-1];
              unloadMuxOut[5] = fifoOut[41][5][w-1];
              unloadMuxOut[6] = fifoOut[42][5][w-1];
              unloadMuxOut[7] = fifoOut[43][5][w-1];
              unloadMuxOut[8] = fifoOut[44][5][w-1];
              unloadMuxOut[9] = fifoOut[45][5][w-1];
              unloadMuxOut[10] = fifoOut[46][5][w-1];
              unloadMuxOut[11] = fifoOut[47][5][w-1];
              unloadMuxOut[12] = fifoOut[48][5][w-1];
              unloadMuxOut[13] = fifoOut[49][5][w-1];
              unloadMuxOut[14] = fifoOut[50][5][w-1];
              unloadMuxOut[15] = fifoOut[51][5][w-1];
              unloadMuxOut[16] = fifoOut[26][4][w-1];
              unloadMuxOut[17] = fifoOut[27][4][w-1];
              unloadMuxOut[18] = fifoOut[28][4][w-1];
              unloadMuxOut[19] = fifoOut[29][4][w-1];
              unloadMuxOut[20] = fifoOut[30][4][w-1];
              unloadMuxOut[21] = fifoOut[31][4][w-1];
              unloadMuxOut[22] = fifoOut[32][4][w-1];
              unloadMuxOut[23] = fifoOut[33][4][w-1];
              unloadMuxOut[24] = fifoOut[34][4][w-1];
              unloadMuxOut[25] = fifoOut[35][4][w-1];
              unloadMuxOut[26] = fifoOut[36][4][w-1];
              unloadMuxOut[27] = fifoOut[37][4][w-1];
              unloadMuxOut[28] = fifoOut[38][4][w-1];
              unloadMuxOut[29] = fifoOut[39][4][w-1];
              unloadMuxOut[30] = fifoOut[40][4][w-1];
              unloadMuxOut[31] = fifoOut[41][4][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[42][4][w-1];
              unloadMuxOut[1] = fifoOut[43][4][w-1];
              unloadMuxOut[2] = fifoOut[44][4][w-1];
              unloadMuxOut[3] = fifoOut[45][4][w-1];
              unloadMuxOut[4] = fifoOut[46][4][w-1];
              unloadMuxOut[5] = fifoOut[47][4][w-1];
              unloadMuxOut[6] = fifoOut[48][4][w-1];
              unloadMuxOut[7] = fifoOut[49][4][w-1];
              unloadMuxOut[8] = fifoOut[50][4][w-1];
              unloadMuxOut[9] = fifoOut[51][4][w-1];
              unloadMuxOut[10] = fifoOut[26][3][w-1];
              unloadMuxOut[11] = fifoOut[27][3][w-1];
              unloadMuxOut[12] = fifoOut[28][3][w-1];
              unloadMuxOut[13] = fifoOut[29][3][w-1];
              unloadMuxOut[14] = fifoOut[30][3][w-1];
              unloadMuxOut[15] = fifoOut[31][3][w-1];
              unloadMuxOut[16] = fifoOut[32][3][w-1];
              unloadMuxOut[17] = fifoOut[33][3][w-1];
              unloadMuxOut[18] = fifoOut[34][3][w-1];
              unloadMuxOut[19] = fifoOut[35][3][w-1];
              unloadMuxOut[20] = fifoOut[36][3][w-1];
              unloadMuxOut[21] = fifoOut[37][3][w-1];
              unloadMuxOut[22] = fifoOut[38][3][w-1];
              unloadMuxOut[23] = fifoOut[39][3][w-1];
              unloadMuxOut[24] = fifoOut[40][3][w-1];
              unloadMuxOut[25] = fifoOut[41][3][w-1];
              unloadMuxOut[26] = fifoOut[42][3][w-1];
              unloadMuxOut[27] = fifoOut[43][3][w-1];
              unloadMuxOut[28] = fifoOut[44][3][w-1];
              unloadMuxOut[29] = fifoOut[45][3][w-1];
              unloadMuxOut[30] = fifoOut[46][3][w-1];
              unloadMuxOut[31] = fifoOut[47][3][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[48][3][w-1];
              unloadMuxOut[1] = fifoOut[49][3][w-1];
              unloadMuxOut[2] = fifoOut[50][3][w-1];
              unloadMuxOut[3] = fifoOut[51][3][w-1];
              unloadMuxOut[4] = fifoOut[26][2][w-1];
              unloadMuxOut[5] = fifoOut[27][2][w-1];
              unloadMuxOut[6] = fifoOut[28][2][w-1];
              unloadMuxOut[7] = fifoOut[29][2][w-1];
              unloadMuxOut[8] = fifoOut[30][2][w-1];
              unloadMuxOut[9] = fifoOut[31][2][w-1];
              unloadMuxOut[10] = fifoOut[32][2][w-1];
              unloadMuxOut[11] = fifoOut[33][2][w-1];
              unloadMuxOut[12] = fifoOut[34][2][w-1];
              unloadMuxOut[13] = fifoOut[35][2][w-1];
              unloadMuxOut[14] = fifoOut[36][2][w-1];
              unloadMuxOut[15] = fifoOut[37][2][w-1];
              unloadMuxOut[16] = fifoOut[38][2][w-1];
              unloadMuxOut[17] = fifoOut[39][2][w-1];
              unloadMuxOut[18] = fifoOut[40][2][w-1];
              unloadMuxOut[19] = fifoOut[41][2][w-1];
              unloadMuxOut[20] = fifoOut[42][2][w-1];
              unloadMuxOut[21] = fifoOut[43][2][w-1];
              unloadMuxOut[22] = fifoOut[44][2][w-1];
              unloadMuxOut[23] = fifoOut[45][2][w-1];
              unloadMuxOut[24] = fifoOut[46][2][w-1];
              unloadMuxOut[25] = fifoOut[47][2][w-1];
              unloadMuxOut[26] = fifoOut[48][2][w-1];
              unloadMuxOut[27] = fifoOut[49][2][w-1];
              unloadMuxOut[28] = fifoOut[50][2][w-1];
              unloadMuxOut[29] = fifoOut[51][2][w-1];
              unloadMuxOut[30] = fifoOut[26][1][w-1];
              unloadMuxOut[31] = fifoOut[27][1][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[28][1][w-1];
              unloadMuxOut[1] = fifoOut[29][1][w-1];
              unloadMuxOut[2] = fifoOut[30][1][w-1];
              unloadMuxOut[3] = fifoOut[31][1][w-1];
              unloadMuxOut[4] = fifoOut[32][1][w-1];
              unloadMuxOut[5] = fifoOut[33][1][w-1];
              unloadMuxOut[6] = fifoOut[34][1][w-1];
              unloadMuxOut[7] = fifoOut[35][1][w-1];
              unloadMuxOut[8] = fifoOut[36][1][w-1];
              unloadMuxOut[9] = fifoOut[37][1][w-1];
              unloadMuxOut[10] = fifoOut[38][1][w-1];
              unloadMuxOut[11] = fifoOut[39][1][w-1];
              unloadMuxOut[12] = fifoOut[40][1][w-1];
              unloadMuxOut[13] = fifoOut[41][1][w-1];
              unloadMuxOut[14] = fifoOut[42][1][w-1];
              unloadMuxOut[15] = fifoOut[43][1][w-1];
              unloadMuxOut[16] = fifoOut[44][1][w-1];
              unloadMuxOut[17] = fifoOut[45][1][w-1];
              unloadMuxOut[18] = fifoOut[46][1][w-1];
              unloadMuxOut[19] = fifoOut[47][1][w-1];
              unloadMuxOut[20] = fifoOut[48][1][w-1];
              unloadMuxOut[21] = fifoOut[49][1][w-1];
              unloadMuxOut[22] = fifoOut[50][1][w-1];
              unloadMuxOut[23] = fifoOut[51][1][w-1];
              unloadMuxOut[24] = fifoOut[26][0][w-1];
              unloadMuxOut[25] = fifoOut[27][0][w-1];
              unloadMuxOut[26] = fifoOut[28][0][w-1];
              unloadMuxOut[27] = fifoOut[29][0][w-1];
              unloadMuxOut[28] = fifoOut[30][0][w-1];
              unloadMuxOut[29] = fifoOut[31][0][w-1];
              unloadMuxOut[30] = fifoOut[32][0][w-1];
              unloadMuxOut[31] = fifoOut[0][11][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[1][11][w-1];
              unloadMuxOut[1] = fifoOut[2][11][w-1];
              unloadMuxOut[2] = fifoOut[3][11][w-1];
              unloadMuxOut[3] = fifoOut[4][11][w-1];
              unloadMuxOut[4] = fifoOut[5][11][w-1];
              unloadMuxOut[5] = fifoOut[6][11][w-1];
              unloadMuxOut[6] = fifoOut[7][11][w-1];
              unloadMuxOut[7] = fifoOut[8][11][w-1];
              unloadMuxOut[8] = fifoOut[9][11][w-1];
              unloadMuxOut[9] = fifoOut[10][11][w-1];
              unloadMuxOut[10] = fifoOut[11][11][w-1];
              unloadMuxOut[11] = fifoOut[12][11][w-1];
              unloadMuxOut[12] = fifoOut[13][11][w-1];
              unloadMuxOut[13] = fifoOut[14][11][w-1];
              unloadMuxOut[14] = fifoOut[15][11][w-1];
              unloadMuxOut[15] = fifoOut[16][11][w-1];
              unloadMuxOut[16] = fifoOut[17][11][w-1];
              unloadMuxOut[17] = fifoOut[18][11][w-1];
              unloadMuxOut[18] = fifoOut[19][11][w-1];
              unloadMuxOut[19] = fifoOut[20][11][w-1];
              unloadMuxOut[20] = fifoOut[21][11][w-1];
              unloadMuxOut[21] = fifoOut[22][11][w-1];
              unloadMuxOut[22] = fifoOut[23][11][w-1];
              unloadMuxOut[23] = fifoOut[24][11][w-1];
              unloadMuxOut[24] = fifoOut[25][11][w-1];
              unloadMuxOut[25] = fifoOut[0][10][w-1];
              unloadMuxOut[26] = fifoOut[1][10][w-1];
              unloadMuxOut[27] = fifoOut[2][10][w-1];
              unloadMuxOut[28] = fifoOut[3][10][w-1];
              unloadMuxOut[29] = fifoOut[4][10][w-1];
              unloadMuxOut[30] = fifoOut[5][10][w-1];
              unloadMuxOut[31] = fifoOut[6][10][w-1];
       end
       16: begin
              unloadMuxOut[0] = fifoOut[7][10][w-1];
              unloadMuxOut[1] = fifoOut[8][10][w-1];
              unloadMuxOut[2] = fifoOut[9][10][w-1];
              unloadMuxOut[3] = fifoOut[10][10][w-1];
              unloadMuxOut[4] = fifoOut[11][10][w-1];
              unloadMuxOut[5] = fifoOut[12][10][w-1];
              unloadMuxOut[6] = fifoOut[13][10][w-1];
              unloadMuxOut[7] = fifoOut[14][10][w-1];
              unloadMuxOut[8] = fifoOut[15][10][w-1];
              unloadMuxOut[9] = fifoOut[16][10][w-1];
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0;
             end
       end
    endcase
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[15][9];
              muxOutConnector[1] = fifoOut[16][9];
              muxOutConnector[2] = fifoOut[17][9];
              muxOutConnector[3] = fifoOut[18][9];
              muxOutConnector[4] = fifoOut[19][9];
              muxOutConnector[5] = fifoOut[20][9];
              muxOutConnector[6] = fifoOut[21][9];
              muxOutConnector[7] = fifoOut[22][9];
              muxOutConnector[8] = fifoOut[23][9];
              muxOutConnector[9] = fifoOut[24][9];
              muxOutConnector[10] = fifoOut[25][9];
              muxOutConnector[11] = fifoOut[0][8];
              muxOutConnector[12] = fifoOut[1][8];
              muxOutConnector[13] = fifoOut[2][8];
              muxOutConnector[14] = fifoOut[3][8];
              muxOutConnector[15] = fifoOut[4][8];
              muxOutConnector[16] = fifoOut[5][8];
              muxOutConnector[17] = fifoOut[6][8];
              muxOutConnector[18] = fifoOut[7][8];
              muxOutConnector[19] = fifoOut[8][8];
              muxOutConnector[20] = fifoOut[9][8];
              muxOutConnector[21] = fifoOut[10][8];
              muxOutConnector[22] = fifoOut[11][8];
              muxOutConnector[23] = fifoOut[12][8];
              muxOutConnector[24] = fifoOut[13][8];
              muxOutConnector[25] = fifoOut[14][8];
              muxOutConnector[26] = fifoOut[48][2];
              muxOutConnector[27] = fifoOut[49][2];
              muxOutConnector[28] = fifoOut[50][2];
              muxOutConnector[29] = fifoOut[51][2];
              muxOutConnector[30] = fifoOut[26][1];
              muxOutConnector[31] = fifoOut[27][1];
              muxOutConnector[32] = fifoOut[28][1];
              muxOutConnector[33] = fifoOut[29][1];
              muxOutConnector[34] = fifoOut[30][1];
              muxOutConnector[35] = fifoOut[31][1];
              muxOutConnector[36] = fifoOut[32][1];
              muxOutConnector[37] = fifoOut[33][1];
              muxOutConnector[38] = fifoOut[34][1];
              muxOutConnector[39] = fifoOut[35][1];
              muxOutConnector[40] = fifoOut[36][1];
              muxOutConnector[41] = fifoOut[37][1];
              muxOutConnector[42] = fifoOut[38][1];
              muxOutConnector[43] = fifoOut[39][1];
              muxOutConnector[44] = fifoOut[40][1];
              muxOutConnector[45] = fifoOut[41][1];
              muxOutConnector[46] = fifoOut[42][1];
              muxOutConnector[47] = fifoOut[43][1];
              muxOutConnector[48] = fifoOut[44][1];
              muxOutConnector[49] = fifoOut[45][1];
              muxOutConnector[50] = fifoOut[46][1];
              muxOutConnector[51] = fifoOut[47][1];
       end
       1: begin
              muxOutConnector[0] = fifoOut[15][8];
              muxOutConnector[1] = fifoOut[16][8];
              muxOutConnector[2] = fifoOut[17][8];
              muxOutConnector[3] = fifoOut[18][8];
              muxOutConnector[4] = fifoOut[19][8];
              muxOutConnector[5] = fifoOut[20][8];
              muxOutConnector[6] = fifoOut[21][8];
              muxOutConnector[7] = fifoOut[22][8];
              muxOutConnector[8] = fifoOut[23][8];
              muxOutConnector[9] = fifoOut[24][8];
              muxOutConnector[10] = fifoOut[25][8];
              muxOutConnector[11] = fifoOut[0][7];
              muxOutConnector[12] = fifoOut[1][7];
              muxOutConnector[13] = fifoOut[2][7];
              muxOutConnector[14] = fifoOut[3][7];
              muxOutConnector[15] = fifoOut[4][7];
              muxOutConnector[16] = fifoOut[5][7];
              muxOutConnector[17] = fifoOut[6][7];
              muxOutConnector[18] = fifoOut[7][7];
              muxOutConnector[19] = fifoOut[8][7];
              muxOutConnector[20] = fifoOut[9][7];
              muxOutConnector[21] = fifoOut[10][7];
              muxOutConnector[22] = fifoOut[11][7];
              muxOutConnector[23] = fifoOut[12][7];
              muxOutConnector[24] = fifoOut[13][7];
              muxOutConnector[25] = fifoOut[14][7];
              muxOutConnector[26] = fifoOut[48][1];
              muxOutConnector[27] = fifoOut[49][1];
              muxOutConnector[28] = fifoOut[50][1];
              muxOutConnector[29] = fifoOut[51][1];
              muxOutConnector[30] = fifoOut[26][0];
              muxOutConnector[31] = fifoOut[27][0];
              muxOutConnector[32] = fifoOut[28][0];
              muxOutConnector[33] = fifoOut[29][0];
              muxOutConnector[34] = fifoOut[30][0];
              muxOutConnector[35] = fifoOut[31][0];
              muxOutConnector[36] = fifoOut[32][0];
              muxOutConnector[37] = fifoOut[0][11];
              muxOutConnector[38] = fifoOut[1][11];
              muxOutConnector[39] = fifoOut[2][11];
              muxOutConnector[40] = fifoOut[3][11];
              muxOutConnector[41] = fifoOut[4][11];
              muxOutConnector[42] = fifoOut[5][11];
              muxOutConnector[43] = fifoOut[6][11];
              muxOutConnector[44] = fifoOut[7][11];
              muxOutConnector[45] = fifoOut[8][11];
              muxOutConnector[46] = fifoOut[9][11];
              muxOutConnector[47] = fifoOut[10][11];
              muxOutConnector[48] = fifoOut[11][11];
              muxOutConnector[49] = fifoOut[12][11];
              muxOutConnector[50] = fifoOut[13][11];
              muxOutConnector[51] = fifoOut[14][11];
       end
       2: begin
              muxOutConnector[0] = fifoOut[15][7];
              muxOutConnector[1] = fifoOut[16][7];
              muxOutConnector[2] = fifoOut[17][7];
              muxOutConnector[3] = fifoOut[18][7];
              muxOutConnector[4] = fifoOut[19][7];
              muxOutConnector[5] = fifoOut[20][7];
              muxOutConnector[6] = fifoOut[21][7];
              muxOutConnector[7] = fifoOut[22][7];
              muxOutConnector[8] = fifoOut[23][7];
              muxOutConnector[9] = fifoOut[24][7];
              muxOutConnector[10] = fifoOut[25][7];
              muxOutConnector[11] = fifoOut[0][6];
              muxOutConnector[12] = fifoOut[1][6];
              muxOutConnector[13] = fifoOut[2][6];
              muxOutConnector[14] = fifoOut[3][6];
              muxOutConnector[15] = fifoOut[4][6];
              muxOutConnector[16] = fifoOut[5][6];
              muxOutConnector[17] = fifoOut[6][6];
              muxOutConnector[18] = fifoOut[7][6];
              muxOutConnector[19] = fifoOut[8][6];
              muxOutConnector[20] = fifoOut[9][6];
              muxOutConnector[21] = fifoOut[10][6];
              muxOutConnector[22] = fifoOut[11][6];
              muxOutConnector[23] = fifoOut[12][6];
              muxOutConnector[24] = fifoOut[13][6];
              muxOutConnector[25] = fifoOut[14][6];
              muxOutConnector[26] = fifoOut[15][11];
              muxOutConnector[27] = fifoOut[16][11];
              muxOutConnector[28] = fifoOut[17][11];
              muxOutConnector[29] = fifoOut[18][11];
              muxOutConnector[30] = fifoOut[19][11];
              muxOutConnector[31] = fifoOut[20][11];
              muxOutConnector[32] = fifoOut[21][11];
              muxOutConnector[33] = fifoOut[22][11];
              muxOutConnector[34] = fifoOut[23][11];
              muxOutConnector[35] = fifoOut[24][11];
              muxOutConnector[36] = fifoOut[25][11];
              muxOutConnector[37] = fifoOut[0][10];
              muxOutConnector[38] = fifoOut[1][10];
              muxOutConnector[39] = fifoOut[2][10];
              muxOutConnector[40] = fifoOut[3][10];
              muxOutConnector[41] = fifoOut[4][10];
              muxOutConnector[42] = fifoOut[5][10];
              muxOutConnector[43] = fifoOut[6][10];
              muxOutConnector[44] = fifoOut[7][10];
              muxOutConnector[45] = fifoOut[8][10];
              muxOutConnector[46] = fifoOut[9][10];
              muxOutConnector[47] = fifoOut[10][10];
              muxOutConnector[48] = fifoOut[11][10];
              muxOutConnector[49] = fifoOut[12][10];
              muxOutConnector[50] = fifoOut[13][10];
              muxOutConnector[51] = fifoOut[14][10];
       end
       3: begin
              muxOutConnector[0] = fifoOut[15][6];
              muxOutConnector[1] = fifoOut[16][6];
              muxOutConnector[2] = fifoOut[17][6];
              muxOutConnector[3] = fifoOut[18][6];
              muxOutConnector[4] = fifoOut[19][6];
              muxOutConnector[5] = fifoOut[20][6];
              muxOutConnector[6] = fifoOut[21][6];
              muxOutConnector[7] = fifoOut[22][6];
              muxOutConnector[8] = fifoOut[23][6];
              muxOutConnector[9] = fifoOut[24][6];
              muxOutConnector[10] = fifoOut[25][6];
              muxOutConnector[11] = fifoOut[0][5];
              muxOutConnector[12] = fifoOut[1][5];
              muxOutConnector[13] = fifoOut[2][5];
              muxOutConnector[14] = fifoOut[3][5];
              muxOutConnector[15] = fifoOut[4][5];
              muxOutConnector[16] = fifoOut[5][5];
              muxOutConnector[17] = fifoOut[6][5];
              muxOutConnector[18] = fifoOut[7][5];
              muxOutConnector[19] = fifoOut[8][5];
              muxOutConnector[20] = fifoOut[9][5];
              muxOutConnector[21] = fifoOut[10][5];
              muxOutConnector[22] = fifoOut[11][5];
              muxOutConnector[23] = fifoOut[12][5];
              muxOutConnector[24] = fifoOut[13][5];
              muxOutConnector[25] = fifoOut[14][5];
              muxOutConnector[26] = fifoOut[15][10];
              muxOutConnector[27] = fifoOut[16][10];
              muxOutConnector[28] = fifoOut[17][10];
              muxOutConnector[29] = fifoOut[18][10];
              muxOutConnector[30] = fifoOut[19][10];
              muxOutConnector[31] = fifoOut[20][10];
              muxOutConnector[32] = fifoOut[21][10];
              muxOutConnector[33] = fifoOut[22][10];
              muxOutConnector[34] = fifoOut[23][10];
              muxOutConnector[35] = fifoOut[24][10];
              muxOutConnector[36] = fifoOut[25][10];
              muxOutConnector[37] = fifoOut[0][9];
              muxOutConnector[38] = fifoOut[1][9];
              muxOutConnector[39] = fifoOut[2][9];
              muxOutConnector[40] = fifoOut[3][9];
              muxOutConnector[41] = fifoOut[4][9];
              muxOutConnector[42] = fifoOut[5][9];
              muxOutConnector[43] = fifoOut[6][9];
              muxOutConnector[44] = fifoOut[7][9];
              muxOutConnector[45] = fifoOut[8][9];
              muxOutConnector[46] = fifoOut[9][9];
              muxOutConnector[47] = fifoOut[10][9];
              muxOutConnector[48] = fifoOut[11][9];
              muxOutConnector[49] = fifoOut[12][9];
              muxOutConnector[50] = fifoOut[13][9];
              muxOutConnector[51] = fifoOut[14][9];
       end
       4: begin
              muxOutConnector[0] = fifoOut[15][5];
              muxOutConnector[1] = fifoOut[16][5];
              muxOutConnector[2] = fifoOut[17][5];
              muxOutConnector[3] = fifoOut[18][5];
              muxOutConnector[4] = fifoOut[19][5];
              muxOutConnector[5] = fifoOut[20][5];
              muxOutConnector[6] = fifoOut[21][5];
              muxOutConnector[7] = fifoOut[22][5];
              muxOutConnector[8] = fifoOut[23][5];
              muxOutConnector[9] = fifoOut[24][5];
              muxOutConnector[10] = fifoOut[25][5];
              muxOutConnector[11] = fifoOut[0][4];
              muxOutConnector[12] = fifoOut[1][4];
              muxOutConnector[13] = fifoOut[2][4];
              muxOutConnector[14] = fifoOut[3][4];
              muxOutConnector[15] = fifoOut[4][4];
              muxOutConnector[16] = fifoOut[5][4];
              muxOutConnector[17] = fifoOut[6][4];
              muxOutConnector[18] = fifoOut[7][4];
              muxOutConnector[19] = fifoOut[8][4];
              muxOutConnector[20] = fifoOut[9][4];
              muxOutConnector[21] = fifoOut[10][4];
              muxOutConnector[22] = fifoOut[11][4];
              muxOutConnector[23] = fifoOut[12][4];
              muxOutConnector[24] = fifoOut[13][4];
              muxOutConnector[25] = fifoOut[14][4];
              muxOutConnector[26] = fifoOut[15][9];
              muxOutConnector[27] = fifoOut[16][9];
              muxOutConnector[28] = fifoOut[17][9];
              muxOutConnector[29] = fifoOut[18][9];
              muxOutConnector[30] = fifoOut[19][9];
              muxOutConnector[31] = fifoOut[20][9];
              muxOutConnector[32] = fifoOut[21][9];
              muxOutConnector[33] = fifoOut[22][9];
              muxOutConnector[34] = fifoOut[23][9];
              muxOutConnector[35] = fifoOut[24][9];
              muxOutConnector[36] = fifoOut[25][9];
              muxOutConnector[37] = fifoOut[0][8];
              muxOutConnector[38] = fifoOut[1][8];
              muxOutConnector[39] = fifoOut[2][8];
              muxOutConnector[40] = fifoOut[3][8];
              muxOutConnector[41] = fifoOut[4][8];
              muxOutConnector[42] = fifoOut[5][8];
              muxOutConnector[43] = fifoOut[6][8];
              muxOutConnector[44] = fifoOut[7][8];
              muxOutConnector[45] = fifoOut[8][8];
              muxOutConnector[46] = fifoOut[9][8];
              muxOutConnector[47] = fifoOut[10][8];
              muxOutConnector[48] = fifoOut[11][8];
              muxOutConnector[49] = fifoOut[12][8];
              muxOutConnector[50] = fifoOut[13][8];
              muxOutConnector[51] = fifoOut[14][8];
       end
       5: begin
              muxOutConnector[0] = fifoOut[15][4];
              muxOutConnector[1] = fifoOut[16][4];
              muxOutConnector[2] = fifoOut[17][4];
              muxOutConnector[3] = fifoOut[18][4];
              muxOutConnector[4] = fifoOut[19][4];
              muxOutConnector[5] = fifoOut[20][4];
              muxOutConnector[6] = fifoOut[21][4];
              muxOutConnector[7] = fifoOut[22][4];
              muxOutConnector[8] = fifoOut[23][4];
              muxOutConnector[9] = fifoOut[24][4];
              muxOutConnector[10] = fifoOut[25][4];
              muxOutConnector[11] = fifoOut[0][3];
              muxOutConnector[12] = fifoOut[1][3];
              muxOutConnector[13] = fifoOut[2][3];
              muxOutConnector[14] = fifoOut[3][3];
              muxOutConnector[15] = fifoOut[4][3];
              muxOutConnector[16] = fifoOut[5][3];
              muxOutConnector[17] = fifoOut[6][3];
              muxOutConnector[18] = fifoOut[7][3];
              muxOutConnector[19] = fifoOut[8][3];
              muxOutConnector[20] = fifoOut[9][3];
              muxOutConnector[21] = fifoOut[26][11];
              muxOutConnector[22] = fifoOut[27][11];
              muxOutConnector[23] = fifoOut[28][11];
              muxOutConnector[24] = fifoOut[29][11];
              muxOutConnector[25] = fifoOut[30][11];
              muxOutConnector[26] = fifoOut[15][8];
              muxOutConnector[27] = fifoOut[16][8];
              muxOutConnector[28] = fifoOut[17][8];
              muxOutConnector[29] = fifoOut[18][8];
              muxOutConnector[30] = fifoOut[19][8];
              muxOutConnector[31] = fifoOut[20][8];
              muxOutConnector[32] = fifoOut[21][8];
              muxOutConnector[33] = fifoOut[22][8];
              muxOutConnector[34] = fifoOut[23][8];
              muxOutConnector[35] = fifoOut[24][8];
              muxOutConnector[36] = fifoOut[25][8];
              muxOutConnector[37] = fifoOut[0][7];
              muxOutConnector[38] = fifoOut[1][7];
              muxOutConnector[39] = fifoOut[2][7];
              muxOutConnector[40] = fifoOut[3][7];
              muxOutConnector[41] = fifoOut[4][7];
              muxOutConnector[42] = fifoOut[5][7];
              muxOutConnector[43] = fifoOut[6][7];
              muxOutConnector[44] = fifoOut[7][7];
              muxOutConnector[45] = fifoOut[8][7];
              muxOutConnector[46] = fifoOut[9][7];
              muxOutConnector[47] = fifoOut[10][7];
              muxOutConnector[48] = fifoOut[11][7];
              muxOutConnector[49] = fifoOut[12][7];
              muxOutConnector[50] = fifoOut[13][7];
              muxOutConnector[51] = fifoOut[14][7];
       end
       6: begin
              muxOutConnector[0] = fifoOut[31][11];
              muxOutConnector[1] = fifoOut[32][11];
              muxOutConnector[2] = fifoOut[33][11];
              muxOutConnector[3] = fifoOut[34][11];
              muxOutConnector[4] = fifoOut[35][11];
              muxOutConnector[5] = fifoOut[36][11];
              muxOutConnector[6] = fifoOut[37][11];
              muxOutConnector[7] = fifoOut[38][11];
              muxOutConnector[8] = fifoOut[39][11];
              muxOutConnector[9] = fifoOut[40][11];
              muxOutConnector[10] = fifoOut[41][11];
              muxOutConnector[11] = fifoOut[42][11];
              muxOutConnector[12] = fifoOut[43][11];
              muxOutConnector[13] = fifoOut[44][11];
              muxOutConnector[14] = fifoOut[45][11];
              muxOutConnector[15] = fifoOut[46][11];
              muxOutConnector[16] = fifoOut[47][11];
              muxOutConnector[17] = fifoOut[48][11];
              muxOutConnector[18] = fifoOut[49][11];
              muxOutConnector[19] = fifoOut[50][11];
              muxOutConnector[20] = fifoOut[51][11];
              muxOutConnector[21] = fifoOut[26][10];
              muxOutConnector[22] = fifoOut[27][10];
              muxOutConnector[23] = fifoOut[28][10];
              muxOutConnector[24] = fifoOut[29][10];
              muxOutConnector[25] = fifoOut[30][10];
              muxOutConnector[26] = fifoOut[15][7];
              muxOutConnector[27] = fifoOut[16][7];
              muxOutConnector[28] = fifoOut[17][7];
              muxOutConnector[29] = fifoOut[18][7];
              muxOutConnector[30] = fifoOut[19][7];
              muxOutConnector[31] = fifoOut[20][7];
              muxOutConnector[32] = fifoOut[21][7];
              muxOutConnector[33] = fifoOut[22][7];
              muxOutConnector[34] = fifoOut[23][7];
              muxOutConnector[35] = fifoOut[24][7];
              muxOutConnector[36] = fifoOut[25][7];
              muxOutConnector[37] = fifoOut[0][6];
              muxOutConnector[38] = fifoOut[1][6];
              muxOutConnector[39] = fifoOut[2][6];
              muxOutConnector[40] = fifoOut[3][6];
              muxOutConnector[41] = fifoOut[4][6];
              muxOutConnector[42] = fifoOut[5][6];
              muxOutConnector[43] = fifoOut[6][6];
              muxOutConnector[44] = fifoOut[7][6];
              muxOutConnector[45] = fifoOut[8][6];
              muxOutConnector[46] = fifoOut[9][6];
              muxOutConnector[47] = fifoOut[10][6];
              muxOutConnector[48] = fifoOut[11][6];
              muxOutConnector[49] = fifoOut[12][6];
              muxOutConnector[50] = fifoOut[13][6];
              muxOutConnector[51] = fifoOut[14][6];
       end
       7: begin
              muxOutConnector[0] = fifoOut[31][10];
              muxOutConnector[1] = fifoOut[32][10];
              muxOutConnector[2] = fifoOut[33][10];
              muxOutConnector[3] = fifoOut[34][10];
              muxOutConnector[4] = fifoOut[35][10];
              muxOutConnector[5] = fifoOut[36][10];
              muxOutConnector[6] = fifoOut[37][10];
              muxOutConnector[7] = fifoOut[38][10];
              muxOutConnector[8] = fifoOut[39][10];
              muxOutConnector[9] = fifoOut[40][10];
              muxOutConnector[10] = fifoOut[41][10];
              muxOutConnector[11] = fifoOut[42][10];
              muxOutConnector[12] = fifoOut[43][10];
              muxOutConnector[13] = fifoOut[44][10];
              muxOutConnector[14] = fifoOut[45][10];
              muxOutConnector[15] = fifoOut[46][10];
              muxOutConnector[16] = fifoOut[47][10];
              muxOutConnector[17] = fifoOut[48][10];
              muxOutConnector[18] = fifoOut[49][10];
              muxOutConnector[19] = fifoOut[50][10];
              muxOutConnector[20] = fifoOut[51][10];
              muxOutConnector[21] = fifoOut[26][9];
              muxOutConnector[22] = fifoOut[27][9];
              muxOutConnector[23] = fifoOut[28][9];
              muxOutConnector[24] = fifoOut[29][9];
              muxOutConnector[25] = fifoOut[30][9];
              muxOutConnector[26] = fifoOut[15][6];
              muxOutConnector[27] = fifoOut[16][6];
              muxOutConnector[28] = fifoOut[17][6];
              muxOutConnector[29] = fifoOut[18][6];
              muxOutConnector[30] = fifoOut[19][6];
              muxOutConnector[31] = fifoOut[20][6];
              muxOutConnector[32] = fifoOut[21][6];
              muxOutConnector[33] = fifoOut[22][6];
              muxOutConnector[34] = fifoOut[23][6];
              muxOutConnector[35] = fifoOut[24][6];
              muxOutConnector[36] = fifoOut[25][6];
              muxOutConnector[37] = fifoOut[0][5];
              muxOutConnector[38] = fifoOut[1][5];
              muxOutConnector[39] = fifoOut[2][5];
              muxOutConnector[40] = fifoOut[3][5];
              muxOutConnector[41] = fifoOut[4][5];
              muxOutConnector[42] = fifoOut[5][5];
              muxOutConnector[43] = fifoOut[6][5];
              muxOutConnector[44] = fifoOut[7][5];
              muxOutConnector[45] = fifoOut[8][5];
              muxOutConnector[46] = fifoOut[9][5];
              muxOutConnector[47] = fifoOut[10][5];
              muxOutConnector[48] = fifoOut[11][5];
              muxOutConnector[49] = fifoOut[12][5];
              muxOutConnector[50] = fifoOut[13][5];
              muxOutConnector[51] = fifoOut[14][5];
       end
       8: begin
              muxOutConnector[0] = fifoOut[31][9];
              muxOutConnector[1] = fifoOut[32][9];
              muxOutConnector[2] = fifoOut[33][9];
              muxOutConnector[3] = fifoOut[34][9];
              muxOutConnector[4] = fifoOut[35][9];
              muxOutConnector[5] = fifoOut[36][9];
              muxOutConnector[6] = fifoOut[37][9];
              muxOutConnector[7] = fifoOut[38][9];
              muxOutConnector[8] = fifoOut[39][9];
              muxOutConnector[9] = fifoOut[40][9];
              muxOutConnector[10] = fifoOut[41][9];
              muxOutConnector[11] = fifoOut[42][9];
              muxOutConnector[12] = fifoOut[43][9];
              muxOutConnector[13] = fifoOut[44][9];
              muxOutConnector[14] = fifoOut[45][9];
              muxOutConnector[15] = fifoOut[46][9];
              muxOutConnector[16] = fifoOut[47][9];
              muxOutConnector[17] = fifoOut[48][9];
              muxOutConnector[18] = fifoOut[49][9];
              muxOutConnector[19] = fifoOut[50][9];
              muxOutConnector[20] = fifoOut[51][9];
              muxOutConnector[21] = fifoOut[26][8];
              muxOutConnector[22] = fifoOut[27][8];
              muxOutConnector[23] = fifoOut[28][8];
              muxOutConnector[24] = fifoOut[29][8];
              muxOutConnector[25] = fifoOut[30][8];
              muxOutConnector[26] = fifoOut[15][5];
              muxOutConnector[27] = fifoOut[16][5];
              muxOutConnector[28] = fifoOut[17][5];
              muxOutConnector[29] = fifoOut[18][5];
              muxOutConnector[30] = fifoOut[19][5];
              muxOutConnector[31] = fifoOut[20][5];
              muxOutConnector[32] = fifoOut[21][5];
              muxOutConnector[33] = fifoOut[22][5];
              muxOutConnector[34] = fifoOut[23][5];
              muxOutConnector[35] = fifoOut[24][5];
              muxOutConnector[36] = fifoOut[25][5];
              muxOutConnector[37] = fifoOut[0][4];
              muxOutConnector[38] = fifoOut[1][4];
              muxOutConnector[39] = fifoOut[2][4];
              muxOutConnector[40] = fifoOut[3][4];
              muxOutConnector[41] = fifoOut[4][4];
              muxOutConnector[42] = fifoOut[5][4];
              muxOutConnector[43] = fifoOut[6][4];
              muxOutConnector[44] = fifoOut[7][4];
              muxOutConnector[45] = fifoOut[8][4];
              muxOutConnector[46] = fifoOut[9][4];
              muxOutConnector[47] = fifoOut[10][4];
              muxOutConnector[48] = fifoOut[11][4];
              muxOutConnector[49] = fifoOut[12][4];
              muxOutConnector[50] = fifoOut[13][4];
              muxOutConnector[51] = fifoOut[14][4];
       end
       9: begin
              muxOutConnector[0] = fifoOut[31][8];
              muxOutConnector[1] = fifoOut[32][8];
              muxOutConnector[2] = fifoOut[33][8];
              muxOutConnector[3] = fifoOut[34][8];
              muxOutConnector[4] = fifoOut[35][8];
              muxOutConnector[5] = fifoOut[36][8];
              muxOutConnector[6] = fifoOut[37][8];
              muxOutConnector[7] = fifoOut[38][8];
              muxOutConnector[8] = fifoOut[39][8];
              muxOutConnector[9] = fifoOut[40][8];
              muxOutConnector[10] = fifoOut[41][8];
              muxOutConnector[11] = fifoOut[42][8];
              muxOutConnector[12] = fifoOut[43][8];
              muxOutConnector[13] = fifoOut[44][8];
              muxOutConnector[14] = fifoOut[45][8];
              muxOutConnector[15] = fifoOut[46][8];
              muxOutConnector[16] = fifoOut[47][8];
              muxOutConnector[17] = fifoOut[48][8];
              muxOutConnector[18] = fifoOut[49][8];
              muxOutConnector[19] = fifoOut[50][8];
              muxOutConnector[20] = fifoOut[51][8];
              muxOutConnector[21] = fifoOut[26][7];
              muxOutConnector[22] = fifoOut[27][7];
              muxOutConnector[23] = fifoOut[28][7];
              muxOutConnector[24] = fifoOut[29][7];
              muxOutConnector[25] = fifoOut[30][7];
              muxOutConnector[26] = fifoOut[15][4];
              muxOutConnector[27] = fifoOut[16][4];
              muxOutConnector[28] = fifoOut[17][4];
              muxOutConnector[29] = fifoOut[18][4];
              muxOutConnector[30] = fifoOut[19][4];
              muxOutConnector[31] = fifoOut[20][4];
              muxOutConnector[32] = fifoOut[21][4];
              muxOutConnector[33] = fifoOut[22][4];
              muxOutConnector[34] = fifoOut[23][4];
              muxOutConnector[35] = fifoOut[24][4];
              muxOutConnector[36] = fifoOut[25][4];
              muxOutConnector[37] = fifoOut[0][3];
              muxOutConnector[38] = fifoOut[1][3];
              muxOutConnector[39] = fifoOut[2][3];
              muxOutConnector[40] = fifoOut[3][3];
              muxOutConnector[41] = fifoOut[4][3];
              muxOutConnector[42] = fifoOut[5][3];
              muxOutConnector[43] = fifoOut[6][3];
              muxOutConnector[44] = fifoOut[7][3];
              muxOutConnector[45] = fifoOut[8][3];
              muxOutConnector[46] = fifoOut[9][3];
              muxOutConnector[47] = fifoOut[26][11];
              muxOutConnector[48] = fifoOut[27][11];
              muxOutConnector[49] = fifoOut[28][11];
              muxOutConnector[50] = fifoOut[29][11];
              muxOutConnector[51] = fifoOut[30][11];
       end
       10: begin
              muxOutConnector[0] = fifoOut[31][7];
              muxOutConnector[1] = fifoOut[32][7];
              muxOutConnector[2] = fifoOut[33][7];
              muxOutConnector[3] = fifoOut[34][7];
              muxOutConnector[4] = fifoOut[35][7];
              muxOutConnector[5] = fifoOut[36][7];
              muxOutConnector[6] = fifoOut[37][7];
              muxOutConnector[7] = fifoOut[38][7];
              muxOutConnector[8] = fifoOut[39][7];
              muxOutConnector[9] = fifoOut[40][7];
              muxOutConnector[10] = fifoOut[41][7];
              muxOutConnector[11] = fifoOut[42][7];
              muxOutConnector[12] = fifoOut[43][7];
              muxOutConnector[13] = fifoOut[44][7];
              muxOutConnector[14] = fifoOut[45][7];
              muxOutConnector[15] = fifoOut[46][7];
              muxOutConnector[16] = fifoOut[47][7];
              muxOutConnector[17] = fifoOut[48][7];
              muxOutConnector[18] = fifoOut[49][7];
              muxOutConnector[19] = fifoOut[50][7];
              muxOutConnector[20] = fifoOut[51][7];
              muxOutConnector[21] = fifoOut[26][6];
              muxOutConnector[22] = fifoOut[27][6];
              muxOutConnector[23] = fifoOut[28][6];
              muxOutConnector[24] = fifoOut[29][6];
              muxOutConnector[25] = fifoOut[30][6];
              muxOutConnector[26] = fifoOut[31][11];
              muxOutConnector[27] = fifoOut[32][11];
              muxOutConnector[28] = fifoOut[33][11];
              muxOutConnector[29] = fifoOut[34][11];
              muxOutConnector[30] = fifoOut[35][11];
              muxOutConnector[31] = fifoOut[36][11];
              muxOutConnector[32] = fifoOut[37][11];
              muxOutConnector[33] = fifoOut[38][11];
              muxOutConnector[34] = fifoOut[39][11];
              muxOutConnector[35] = fifoOut[40][11];
              muxOutConnector[36] = fifoOut[41][11];
              muxOutConnector[37] = fifoOut[42][11];
              muxOutConnector[38] = fifoOut[43][11];
              muxOutConnector[39] = fifoOut[44][11];
              muxOutConnector[40] = fifoOut[45][11];
              muxOutConnector[41] = fifoOut[46][11];
              muxOutConnector[42] = fifoOut[47][11];
              muxOutConnector[43] = fifoOut[48][11];
              muxOutConnector[44] = fifoOut[49][11];
              muxOutConnector[45] = fifoOut[50][11];
              muxOutConnector[46] = fifoOut[51][11];
              muxOutConnector[47] = fifoOut[26][10];
              muxOutConnector[48] = fifoOut[27][10];
              muxOutConnector[49] = fifoOut[28][10];
              muxOutConnector[50] = fifoOut[29][10];
              muxOutConnector[51] = fifoOut[30][10];
       end
       11: begin
              muxOutConnector[0] = fifoOut[31][6];
              muxOutConnector[1] = fifoOut[32][6];
              muxOutConnector[2] = fifoOut[33][6];
              muxOutConnector[3] = fifoOut[34][6];
              muxOutConnector[4] = fifoOut[35][6];
              muxOutConnector[5] = fifoOut[36][6];
              muxOutConnector[6] = fifoOut[37][6];
              muxOutConnector[7] = fifoOut[38][6];
              muxOutConnector[8] = fifoOut[39][6];
              muxOutConnector[9] = fifoOut[40][6];
              muxOutConnector[10] = fifoOut[41][6];
              muxOutConnector[11] = fifoOut[42][6];
              muxOutConnector[12] = fifoOut[43][6];
              muxOutConnector[13] = fifoOut[44][6];
              muxOutConnector[14] = fifoOut[45][6];
              muxOutConnector[15] = fifoOut[46][6];
              muxOutConnector[16] = fifoOut[47][6];
              muxOutConnector[17] = fifoOut[48][6];
              muxOutConnector[18] = fifoOut[49][6];
              muxOutConnector[19] = fifoOut[50][6];
              muxOutConnector[20] = fifoOut[51][6];
              muxOutConnector[21] = fifoOut[26][5];
              muxOutConnector[22] = fifoOut[27][5];
              muxOutConnector[23] = fifoOut[28][5];
              muxOutConnector[24] = fifoOut[29][5];
              muxOutConnector[25] = fifoOut[30][5];
              muxOutConnector[26] = fifoOut[31][10];
              muxOutConnector[27] = fifoOut[32][10];
              muxOutConnector[28] = fifoOut[33][10];
              muxOutConnector[29] = fifoOut[34][10];
              muxOutConnector[30] = fifoOut[35][10];
              muxOutConnector[31] = fifoOut[36][10];
              muxOutConnector[32] = fifoOut[37][10];
              muxOutConnector[33] = fifoOut[38][10];
              muxOutConnector[34] = fifoOut[39][10];
              muxOutConnector[35] = fifoOut[40][10];
              muxOutConnector[36] = fifoOut[41][10];
              muxOutConnector[37] = fifoOut[42][10];
              muxOutConnector[38] = fifoOut[43][10];
              muxOutConnector[39] = fifoOut[44][10];
              muxOutConnector[40] = fifoOut[45][10];
              muxOutConnector[41] = fifoOut[46][10];
              muxOutConnector[42] = fifoOut[47][10];
              muxOutConnector[43] = fifoOut[48][10];
              muxOutConnector[44] = fifoOut[49][10];
              muxOutConnector[45] = fifoOut[50][10];
              muxOutConnector[46] = fifoOut[51][10];
              muxOutConnector[47] = fifoOut[26][9];
              muxOutConnector[48] = fifoOut[27][9];
              muxOutConnector[49] = fifoOut[28][9];
              muxOutConnector[50] = fifoOut[29][9];
              muxOutConnector[51] = fifoOut[30][9];
       end
       12: begin
              muxOutConnector[0] = fifoOut[31][5];
              muxOutConnector[1] = fifoOut[32][5];
              muxOutConnector[2] = fifoOut[33][5];
              muxOutConnector[3] = fifoOut[34][5];
              muxOutConnector[4] = fifoOut[35][5];
              muxOutConnector[5] = fifoOut[36][5];
              muxOutConnector[6] = fifoOut[37][5];
              muxOutConnector[7] = fifoOut[38][5];
              muxOutConnector[8] = fifoOut[39][5];
              muxOutConnector[9] = fifoOut[40][5];
              muxOutConnector[10] = fifoOut[41][5];
              muxOutConnector[11] = fifoOut[42][5];
              muxOutConnector[12] = fifoOut[43][5];
              muxOutConnector[13] = fifoOut[44][5];
              muxOutConnector[14] = fifoOut[45][5];
              muxOutConnector[15] = fifoOut[46][5];
              muxOutConnector[16] = fifoOut[47][5];
              muxOutConnector[17] = fifoOut[48][5];
              muxOutConnector[18] = fifoOut[49][5];
              muxOutConnector[19] = fifoOut[50][5];
              muxOutConnector[20] = fifoOut[51][5];
              muxOutConnector[21] = fifoOut[26][4];
              muxOutConnector[22] = fifoOut[27][4];
              muxOutConnector[23] = fifoOut[28][4];
              muxOutConnector[24] = fifoOut[29][4];
              muxOutConnector[25] = fifoOut[30][4];
              muxOutConnector[26] = fifoOut[31][9];
              muxOutConnector[27] = fifoOut[32][9];
              muxOutConnector[28] = fifoOut[33][9];
              muxOutConnector[29] = fifoOut[34][9];
              muxOutConnector[30] = fifoOut[35][9];
              muxOutConnector[31] = fifoOut[36][9];
              muxOutConnector[32] = fifoOut[37][9];
              muxOutConnector[33] = fifoOut[38][9];
              muxOutConnector[34] = fifoOut[39][9];
              muxOutConnector[35] = fifoOut[40][9];
              muxOutConnector[36] = fifoOut[41][9];
              muxOutConnector[37] = fifoOut[42][9];
              muxOutConnector[38] = fifoOut[43][9];
              muxOutConnector[39] = fifoOut[44][9];
              muxOutConnector[40] = fifoOut[45][9];
              muxOutConnector[41] = fifoOut[46][9];
              muxOutConnector[42] = fifoOut[47][9];
              muxOutConnector[43] = fifoOut[48][9];
              muxOutConnector[44] = fifoOut[49][9];
              muxOutConnector[45] = fifoOut[50][9];
              muxOutConnector[46] = fifoOut[51][9];
              muxOutConnector[47] = fifoOut[26][8];
              muxOutConnector[48] = fifoOut[27][8];
              muxOutConnector[49] = fifoOut[28][8];
              muxOutConnector[50] = fifoOut[29][8];
              muxOutConnector[51] = fifoOut[30][8];
       end
       13: begin
              muxOutConnector[0] = fifoOut[31][4];
              muxOutConnector[1] = fifoOut[32][4];
              muxOutConnector[2] = fifoOut[33][4];
              muxOutConnector[3] = fifoOut[34][4];
              muxOutConnector[4] = fifoOut[35][4];
              muxOutConnector[5] = fifoOut[36][4];
              muxOutConnector[6] = fifoOut[37][4];
              muxOutConnector[7] = fifoOut[38][4];
              muxOutConnector[8] = fifoOut[39][4];
              muxOutConnector[9] = fifoOut[40][4];
              muxOutConnector[10] = fifoOut[41][4];
              muxOutConnector[11] = fifoOut[42][4];
              muxOutConnector[12] = fifoOut[43][4];
              muxOutConnector[13] = fifoOut[44][4];
              muxOutConnector[14] = fifoOut[45][4];
              muxOutConnector[15] = fifoOut[46][4];
              muxOutConnector[16] = fifoOut[47][4];
              muxOutConnector[17] = fifoOut[48][4];
              muxOutConnector[18] = fifoOut[49][4];
              muxOutConnector[19] = fifoOut[50][4];
              muxOutConnector[20] = fifoOut[51][4];
              muxOutConnector[21] = fifoOut[26][3];
              muxOutConnector[22] = fifoOut[27][3];
              muxOutConnector[23] = fifoOut[28][3];
              muxOutConnector[24] = fifoOut[29][3];
              muxOutConnector[25] = fifoOut[30][3];
              muxOutConnector[26] = fifoOut[31][8];
              muxOutConnector[27] = fifoOut[32][8];
              muxOutConnector[28] = fifoOut[33][8];
              muxOutConnector[29] = fifoOut[34][8];
              muxOutConnector[30] = fifoOut[35][8];
              muxOutConnector[31] = fifoOut[36][8];
              muxOutConnector[32] = fifoOut[37][8];
              muxOutConnector[33] = fifoOut[38][8];
              muxOutConnector[34] = fifoOut[39][8];
              muxOutConnector[35] = fifoOut[40][8];
              muxOutConnector[36] = fifoOut[41][8];
              muxOutConnector[37] = fifoOut[42][8];
              muxOutConnector[38] = fifoOut[43][8];
              muxOutConnector[39] = fifoOut[44][8];
              muxOutConnector[40] = fifoOut[45][8];
              muxOutConnector[41] = fifoOut[46][8];
              muxOutConnector[42] = fifoOut[47][8];
              muxOutConnector[43] = fifoOut[48][8];
              muxOutConnector[44] = fifoOut[49][8];
              muxOutConnector[45] = fifoOut[50][8];
              muxOutConnector[46] = fifoOut[51][8];
              muxOutConnector[47] = fifoOut[26][7];
              muxOutConnector[48] = fifoOut[27][7];
              muxOutConnector[49] = fifoOut[28][7];
              muxOutConnector[50] = fifoOut[29][7];
              muxOutConnector[51] = fifoOut[30][7];
       end
       14: begin
              muxOutConnector[0] = fifoOut[31][3];
              muxOutConnector[1] = fifoOut[32][3];
              muxOutConnector[2] = fifoOut[33][3];
              muxOutConnector[3] = fifoOut[34][3];
              muxOutConnector[4] = fifoOut[35][3];
              muxOutConnector[5] = fifoOut[36][3];
              muxOutConnector[6] = fifoOut[37][3];
              muxOutConnector[7] = fifoOut[38][3];
              muxOutConnector[8] = fifoOut[39][3];
              muxOutConnector[9] = fifoOut[40][3];
              muxOutConnector[10] = fifoOut[41][3];
              muxOutConnector[11] = fifoOut[42][3];
              muxOutConnector[12] = fifoOut[43][3];
              muxOutConnector[13] = fifoOut[44][3];
              muxOutConnector[14] = fifoOut[45][3];
              muxOutConnector[15] = fifoOut[46][3];
              muxOutConnector[16] = fifoOut[47][3];
              muxOutConnector[17] = fifoOut[48][3];
              muxOutConnector[18] = fifoOut[49][3];
              muxOutConnector[19] = fifoOut[50][3];
              muxOutConnector[20] = fifoOut[51][3];
              muxOutConnector[21] = fifoOut[26][2];
              muxOutConnector[22] = fifoOut[27][2];
              muxOutConnector[23] = fifoOut[28][2];
              muxOutConnector[24] = fifoOut[29][2];
              muxOutConnector[25] = fifoOut[30][2];
              muxOutConnector[26] = fifoOut[31][7];
              muxOutConnector[27] = fifoOut[32][7];
              muxOutConnector[28] = fifoOut[33][7];
              muxOutConnector[29] = fifoOut[34][7];
              muxOutConnector[30] = fifoOut[35][7];
              muxOutConnector[31] = fifoOut[36][7];
              muxOutConnector[32] = fifoOut[37][7];
              muxOutConnector[33] = fifoOut[38][7];
              muxOutConnector[34] = fifoOut[39][7];
              muxOutConnector[35] = fifoOut[40][7];
              muxOutConnector[36] = fifoOut[41][7];
              muxOutConnector[37] = fifoOut[42][7];
              muxOutConnector[38] = fifoOut[43][7];
              muxOutConnector[39] = fifoOut[44][7];
              muxOutConnector[40] = fifoOut[45][7];
              muxOutConnector[41] = fifoOut[46][7];
              muxOutConnector[42] = fifoOut[47][7];
              muxOutConnector[43] = fifoOut[48][7];
              muxOutConnector[44] = fifoOut[49][7];
              muxOutConnector[45] = fifoOut[50][7];
              muxOutConnector[46] = fifoOut[51][7];
              muxOutConnector[47] = fifoOut[26][6];
              muxOutConnector[48] = fifoOut[27][6];
              muxOutConnector[49] = fifoOut[28][6];
              muxOutConnector[50] = fifoOut[29][6];
              muxOutConnector[51] = fifoOut[30][6];
       end
       15: begin
              muxOutConnector[0] = fifoOut[31][2];
              muxOutConnector[1] = fifoOut[32][2];
              muxOutConnector[2] = fifoOut[33][2];
              muxOutConnector[3] = fifoOut[34][2];
              muxOutConnector[4] = fifoOut[35][2];
              muxOutConnector[5] = fifoOut[36][2];
              muxOutConnector[6] = fifoOut[37][2];
              muxOutConnector[7] = fifoOut[38][2];
              muxOutConnector[8] = fifoOut[39][2];
              muxOutConnector[9] = fifoOut[40][2];
              muxOutConnector[10] = fifoOut[41][2];
              muxOutConnector[11] = fifoOut[42][2];
              muxOutConnector[12] = fifoOut[43][2];
              muxOutConnector[13] = fifoOut[44][2];
              muxOutConnector[14] = fifoOut[45][2];
              muxOutConnector[15] = fifoOut[46][2];
              muxOutConnector[16] = fifoOut[47][2];
              muxOutConnector[17] = fifoOut[48][2];
              muxOutConnector[18] = fifoOut[49][2];
              muxOutConnector[19] = fifoOut[50][2];
              muxOutConnector[20] = fifoOut[51][2];
              muxOutConnector[21] = fifoOut[26][1];
              muxOutConnector[22] = fifoOut[27][1];
              muxOutConnector[23] = fifoOut[28][1];
              muxOutConnector[24] = fifoOut[29][1];
              muxOutConnector[25] = fifoOut[30][1];
              muxOutConnector[26] = fifoOut[31][6];
              muxOutConnector[27] = fifoOut[32][6];
              muxOutConnector[28] = fifoOut[33][6];
              muxOutConnector[29] = fifoOut[34][6];
              muxOutConnector[30] = fifoOut[35][6];
              muxOutConnector[31] = fifoOut[36][6];
              muxOutConnector[32] = fifoOut[37][6];
              muxOutConnector[33] = fifoOut[38][6];
              muxOutConnector[34] = fifoOut[39][6];
              muxOutConnector[35] = fifoOut[40][6];
              muxOutConnector[36] = fifoOut[41][6];
              muxOutConnector[37] = fifoOut[42][6];
              muxOutConnector[38] = fifoOut[43][6];
              muxOutConnector[39] = fifoOut[44][6];
              muxOutConnector[40] = fifoOut[45][6];
              muxOutConnector[41] = fifoOut[46][6];
              muxOutConnector[42] = fifoOut[47][6];
              muxOutConnector[43] = fifoOut[48][6];
              muxOutConnector[44] = fifoOut[49][6];
              muxOutConnector[45] = fifoOut[50][6];
              muxOutConnector[46] = fifoOut[51][6];
              muxOutConnector[47] = fifoOut[26][5];
              muxOutConnector[48] = fifoOut[27][5];
              muxOutConnector[49] = fifoOut[28][5];
              muxOutConnector[50] = fifoOut[29][5];
              muxOutConnector[51] = fifoOut[30][5];
       end
       16: begin
              muxOutConnector[0] = fifoOut[31][1];
              muxOutConnector[1] = fifoOut[32][1];
              muxOutConnector[2] = fifoOut[33][1];
              muxOutConnector[3] = fifoOut[34][1];
              muxOutConnector[4] = fifoOut[35][1];
              muxOutConnector[5] = fifoOut[36][1];
              muxOutConnector[6] = fifoOut[37][1];
              muxOutConnector[7] = fifoOut[38][1];
              muxOutConnector[8] = fifoOut[39][1];
              muxOutConnector[9] = fifoOut[40][1];
              muxOutConnector[10] = fifoOut[41][1];
              muxOutConnector[11] = fifoOut[42][1];
              muxOutConnector[12] = fifoOut[43][1];
              muxOutConnector[13] = fifoOut[44][1];
              muxOutConnector[14] = fifoOut[45][1];
              muxOutConnector[15] = fifoOut[46][1];
              muxOutConnector[16] = fifoOut[47][1];
              muxOutConnector[17] = fifoOut[48][1];
              muxOutConnector[18] = fifoOut[49][1];
              muxOutConnector[19] = fifoOut[50][1];
              muxOutConnector[20] = fifoOut[51][1];
              muxOutConnector[21] = fifoOut[26][0];
              muxOutConnector[22] = fifoOut[27][0];
              muxOutConnector[23] = fifoOut[28][0];
              muxOutConnector[24] = fifoOut[29][0];
              muxOutConnector[25] = fifoOut[30][0];
              muxOutConnector[26] = fifoOut[31][5];
              muxOutConnector[27] = fifoOut[32][5];
              muxOutConnector[28] = fifoOut[33][5];
              muxOutConnector[29] = fifoOut[34][5];
              muxOutConnector[30] = fifoOut[35][5];
              muxOutConnector[31] = fifoOut[36][5];
              muxOutConnector[32] = fifoOut[37][5];
              muxOutConnector[33] = fifoOut[38][5];
              muxOutConnector[34] = fifoOut[39][5];
              muxOutConnector[35] = fifoOut[40][5];
              muxOutConnector[36] = fifoOut[41][5];
              muxOutConnector[37] = fifoOut[42][5];
              muxOutConnector[38] = fifoOut[43][5];
              muxOutConnector[39] = fifoOut[44][5];
              muxOutConnector[40] = fifoOut[45][5];
              muxOutConnector[41] = fifoOut[46][5];
              muxOutConnector[42] = fifoOut[47][5];
              muxOutConnector[43] = fifoOut[48][5];
              muxOutConnector[44] = fifoOut[49][5];
              muxOutConnector[45] = fifoOut[50][5];
              muxOutConnector[46] = fifoOut[51][5];
              muxOutConnector[47] = fifoOut[26][4];
              muxOutConnector[48] = fifoOut[27][4];
              muxOutConnector[49] = fifoOut[28][4];
              muxOutConnector[50] = fifoOut[29][4];
              muxOutConnector[51] = fifoOut[30][4];
       end
       17: begin
              muxOutConnector[0] = fifoOut[31][0];
              muxOutConnector[1] = fifoOut[32][0];
              muxOutConnector[2] = fifoOut[0][11];
              muxOutConnector[3] = fifoOut[1][11];
              muxOutConnector[4] = fifoOut[2][11];
              muxOutConnector[5] = fifoOut[3][11];
              muxOutConnector[6] = fifoOut[4][11];
              muxOutConnector[7] = fifoOut[5][11];
              muxOutConnector[8] = fifoOut[6][11];
              muxOutConnector[9] = fifoOut[7][11];
              muxOutConnector[10] = fifoOut[8][11];
              muxOutConnector[11] = fifoOut[9][11];
              muxOutConnector[12] = fifoOut[10][11];
              muxOutConnector[13] = fifoOut[11][11];
              muxOutConnector[14] = fifoOut[12][11];
              muxOutConnector[15] = fifoOut[13][11];
              muxOutConnector[16] = fifoOut[14][11];
              muxOutConnector[17] = fifoOut[15][11];
              muxOutConnector[18] = fifoOut[16][11];
              muxOutConnector[19] = fifoOut[17][11];
              muxOutConnector[20] = fifoOut[18][11];
              muxOutConnector[21] = fifoOut[19][11];
              muxOutConnector[22] = fifoOut[20][11];
              muxOutConnector[23] = fifoOut[21][11];
              muxOutConnector[24] = fifoOut[22][11];
              muxOutConnector[25] = fifoOut[23][11];
              muxOutConnector[26] = fifoOut[31][4];
              muxOutConnector[27] = fifoOut[32][4];
              muxOutConnector[28] = fifoOut[33][4];
              muxOutConnector[29] = fifoOut[34][4];
              muxOutConnector[30] = fifoOut[35][4];
              muxOutConnector[31] = fifoOut[36][4];
              muxOutConnector[32] = fifoOut[37][4];
              muxOutConnector[33] = fifoOut[38][4];
              muxOutConnector[34] = fifoOut[39][4];
              muxOutConnector[35] = fifoOut[40][4];
              muxOutConnector[36] = fifoOut[41][4];
              muxOutConnector[37] = fifoOut[42][4];
              muxOutConnector[38] = fifoOut[43][4];
              muxOutConnector[39] = fifoOut[44][4];
              muxOutConnector[40] = fifoOut[45][4];
              muxOutConnector[41] = fifoOut[46][4];
              muxOutConnector[42] = fifoOut[47][4];
              muxOutConnector[43] = fifoOut[48][4];
              muxOutConnector[44] = fifoOut[49][4];
              muxOutConnector[45] = fifoOut[50][4];
              muxOutConnector[46] = fifoOut[51][4];
              muxOutConnector[47] = fifoOut[26][3];
              muxOutConnector[48] = fifoOut[27][3];
              muxOutConnector[49] = fifoOut[28][3];
              muxOutConnector[50] = fifoOut[29][3];
              muxOutConnector[51] = fifoOut[30][3];
       end
       18: begin
              muxOutConnector[0] = fifoOut[24][11];
              muxOutConnector[1] = fifoOut[25][11];
              muxOutConnector[2] = fifoOut[0][10];
              muxOutConnector[3] = fifoOut[1][10];
              muxOutConnector[4] = fifoOut[2][10];
              muxOutConnector[5] = fifoOut[3][10];
              muxOutConnector[6] = fifoOut[4][10];
              muxOutConnector[7] = fifoOut[5][10];
              muxOutConnector[8] = fifoOut[6][10];
              muxOutConnector[9] = fifoOut[7][10];
              muxOutConnector[10] = fifoOut[8][10];
              muxOutConnector[11] = fifoOut[9][10];
              muxOutConnector[12] = fifoOut[10][10];
              muxOutConnector[13] = fifoOut[11][10];
              muxOutConnector[14] = fifoOut[12][10];
              muxOutConnector[15] = fifoOut[13][10];
              muxOutConnector[16] = fifoOut[14][10];
              muxOutConnector[17] = fifoOut[15][10];
              muxOutConnector[18] = fifoOut[16][10];
              muxOutConnector[19] = fifoOut[17][10];
              muxOutConnector[20] = fifoOut[18][10];
              muxOutConnector[21] = fifoOut[19][10];
              muxOutConnector[22] = fifoOut[20][10];
              muxOutConnector[23] = fifoOut[21][10];
              muxOutConnector[24] = fifoOut[22][10];
              muxOutConnector[25] = fifoOut[23][10];
              muxOutConnector[26] = fifoOut[31][3];
              muxOutConnector[27] = fifoOut[32][3];
              muxOutConnector[28] = fifoOut[33][3];
              muxOutConnector[29] = fifoOut[34][3];
              muxOutConnector[30] = fifoOut[35][3];
              muxOutConnector[31] = fifoOut[36][3];
              muxOutConnector[32] = fifoOut[37][3];
              muxOutConnector[33] = fifoOut[38][3];
              muxOutConnector[34] = fifoOut[39][3];
              muxOutConnector[35] = fifoOut[40][3];
              muxOutConnector[36] = fifoOut[41][3];
              muxOutConnector[37] = fifoOut[42][3];
              muxOutConnector[38] = fifoOut[43][3];
              muxOutConnector[39] = fifoOut[44][3];
              muxOutConnector[40] = fifoOut[45][3];
              muxOutConnector[41] = fifoOut[46][3];
              muxOutConnector[42] = fifoOut[47][3];
              muxOutConnector[43] = fifoOut[48][3];
              muxOutConnector[44] = fifoOut[49][3];
              muxOutConnector[45] = fifoOut[50][3];
              muxOutConnector[46] = fifoOut[51][3];
              muxOutConnector[47] = fifoOut[26][2];
              muxOutConnector[48] = fifoOut[27][2];
              muxOutConnector[49] = fifoOut[28][2];
              muxOutConnector[50] = fifoOut[29][2];
              muxOutConnector[51] = fifoOut[30][2];
       end
       19: begin
              muxOutConnector[0] = fifoOut[24][10];
              muxOutConnector[1] = fifoOut[25][10];
              muxOutConnector[2] = fifoOut[0][9];
              muxOutConnector[3] = fifoOut[1][9];
              muxOutConnector[4] = fifoOut[2][9];
              muxOutConnector[5] = fifoOut[3][9];
              muxOutConnector[6] = fifoOut[4][9];
              muxOutConnector[7] = fifoOut[5][9];
              muxOutConnector[8] = fifoOut[6][9];
              muxOutConnector[9] = fifoOut[7][9];
              muxOutConnector[10] = fifoOut[8][9];
              muxOutConnector[11] = fifoOut[9][9];
              muxOutConnector[12] = fifoOut[10][9];
              muxOutConnector[13] = fifoOut[11][9];
              muxOutConnector[14] = fifoOut[12][9];
              muxOutConnector[15] = fifoOut[13][9];
              muxOutConnector[16] = fifoOut[14][9];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[31][2];
              muxOutConnector[27] = fifoOut[32][2];
              muxOutConnector[28] = fifoOut[33][2];
              muxOutConnector[29] = fifoOut[34][2];
              muxOutConnector[30] = fifoOut[35][2];
              muxOutConnector[31] = fifoOut[36][2];
              muxOutConnector[32] = fifoOut[37][2];
              muxOutConnector[33] = fifoOut[38][2];
              muxOutConnector[34] = fifoOut[39][2];
              muxOutConnector[35] = fifoOut[40][2];
              muxOutConnector[36] = fifoOut[41][2];
              muxOutConnector[37] = fifoOut[42][2];
              muxOutConnector[38] = fifoOut[43][2];
              muxOutConnector[39] = fifoOut[44][2];
              muxOutConnector[40] = fifoOut[45][2];
              muxOutConnector[41] = fifoOut[46][2];
              muxOutConnector[42] = fifoOut[47][2];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
