`timescale 1ns / 1ps
module LMem1To0_511_circ3_yesshift_nounload_scripted(
        muxOut,
        ly0In,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 12;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            fifoOut[i][0] <= ly0InConnector[i];
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[15][9];
              muxOutConnector[1] = fifoOut[16][9];
              muxOutConnector[2] = fifoOut[17][9];
              muxOutConnector[3] = fifoOut[18][9];
              muxOutConnector[4] = fifoOut[19][9];
              muxOutConnector[5] = fifoOut[20][9];
              muxOutConnector[6] = fifoOut[21][9];
              muxOutConnector[7] = fifoOut[22][9];
              muxOutConnector[8] = fifoOut[23][9];
              muxOutConnector[9] = fifoOut[24][9];
              muxOutConnector[10] = fifoOut[25][9];
              muxOutConnector[11] = fifoOut[0][8];
              muxOutConnector[12] = fifoOut[1][8];
              muxOutConnector[13] = fifoOut[2][8];
              muxOutConnector[14] = fifoOut[3][8];
              muxOutConnector[15] = fifoOut[4][8];
              muxOutConnector[16] = fifoOut[5][8];
              muxOutConnector[17] = fifoOut[6][8];
              muxOutConnector[18] = fifoOut[7][8];
              muxOutConnector[19] = fifoOut[8][8];
              muxOutConnector[20] = fifoOut[9][8];
              muxOutConnector[21] = fifoOut[10][8];
              muxOutConnector[22] = fifoOut[11][8];
              muxOutConnector[23] = fifoOut[12][8];
              muxOutConnector[24] = fifoOut[13][8];
              muxOutConnector[25] = fifoOut[14][8];
              muxOutConnector[26] = fifoOut[48][2];
              muxOutConnector[27] = fifoOut[49][2];
              muxOutConnector[28] = fifoOut[50][2];
              muxOutConnector[29] = fifoOut[51][2];
              muxOutConnector[30] = fifoOut[26][1];
              muxOutConnector[31] = fifoOut[27][1];
              muxOutConnector[32] = fifoOut[28][1];
              muxOutConnector[33] = fifoOut[29][1];
              muxOutConnector[34] = fifoOut[30][1];
              muxOutConnector[35] = fifoOut[31][1];
              muxOutConnector[36] = fifoOut[32][1];
              muxOutConnector[37] = fifoOut[33][1];
              muxOutConnector[38] = fifoOut[34][1];
              muxOutConnector[39] = fifoOut[35][1];
              muxOutConnector[40] = fifoOut[36][1];
              muxOutConnector[41] = fifoOut[37][1];
              muxOutConnector[42] = fifoOut[38][1];
              muxOutConnector[43] = fifoOut[39][1];
              muxOutConnector[44] = fifoOut[40][1];
              muxOutConnector[45] = fifoOut[41][1];
              muxOutConnector[46] = fifoOut[42][1];
              muxOutConnector[47] = fifoOut[43][1];
              muxOutConnector[48] = fifoOut[44][1];
              muxOutConnector[49] = fifoOut[45][1];
              muxOutConnector[50] = fifoOut[46][1];
              muxOutConnector[51] = fifoOut[47][1];
       end
       1: begin
              muxOutConnector[0] = fifoOut[15][9];
              muxOutConnector[1] = fifoOut[16][9];
              muxOutConnector[2] = fifoOut[17][9];
              muxOutConnector[3] = fifoOut[18][9];
              muxOutConnector[4] = fifoOut[19][9];
              muxOutConnector[5] = fifoOut[20][9];
              muxOutConnector[6] = fifoOut[21][9];
              muxOutConnector[7] = fifoOut[22][9];
              muxOutConnector[8] = fifoOut[23][9];
              muxOutConnector[9] = fifoOut[24][9];
              muxOutConnector[10] = fifoOut[25][9];
              muxOutConnector[11] = fifoOut[0][8];
              muxOutConnector[12] = fifoOut[1][8];
              muxOutConnector[13] = fifoOut[2][8];
              muxOutConnector[14] = fifoOut[3][8];
              muxOutConnector[15] = fifoOut[4][8];
              muxOutConnector[16] = fifoOut[5][8];
              muxOutConnector[17] = fifoOut[6][8];
              muxOutConnector[18] = fifoOut[7][8];
              muxOutConnector[19] = fifoOut[8][8];
              muxOutConnector[20] = fifoOut[9][8];
              muxOutConnector[21] = fifoOut[10][8];
              muxOutConnector[22] = fifoOut[11][8];
              muxOutConnector[23] = fifoOut[12][8];
              muxOutConnector[24] = fifoOut[13][8];
              muxOutConnector[25] = fifoOut[14][8];
              muxOutConnector[26] = fifoOut[48][2];
              muxOutConnector[27] = fifoOut[49][2];
              muxOutConnector[28] = fifoOut[50][2];
              muxOutConnector[29] = fifoOut[51][2];
              muxOutConnector[30] = fifoOut[26][1];
              muxOutConnector[31] = fifoOut[27][1];
              muxOutConnector[32] = fifoOut[28][1];
              muxOutConnector[33] = fifoOut[29][1];
              muxOutConnector[34] = fifoOut[30][1];
              muxOutConnector[35] = fifoOut[31][1];
              muxOutConnector[36] = fifoOut[32][1];
              muxOutConnector[37] = fifoOut[33][1];
              muxOutConnector[38] = fifoOut[34][1];
              muxOutConnector[39] = fifoOut[35][1];
              muxOutConnector[40] = fifoOut[36][1];
              muxOutConnector[41] = fifoOut[37][1];
              muxOutConnector[42] = fifoOut[38][1];
              muxOutConnector[43] = fifoOut[39][1];
              muxOutConnector[44] = fifoOut[40][1];
              muxOutConnector[45] = fifoOut[41][1];
              muxOutConnector[46] = fifoOut[42][1];
              muxOutConnector[47] = fifoOut[10][0];
              muxOutConnector[48] = fifoOut[11][0];
              muxOutConnector[49] = fifoOut[12][0];
              muxOutConnector[50] = fifoOut[13][0];
              muxOutConnector[51] = fifoOut[14][0];
       end
       2: begin
              muxOutConnector[0] = fifoOut[15][9];
              muxOutConnector[1] = fifoOut[16][9];
              muxOutConnector[2] = fifoOut[17][9];
              muxOutConnector[3] = fifoOut[18][9];
              muxOutConnector[4] = fifoOut[19][9];
              muxOutConnector[5] = fifoOut[20][9];
              muxOutConnector[6] = fifoOut[21][9];
              muxOutConnector[7] = fifoOut[22][9];
              muxOutConnector[8] = fifoOut[23][9];
              muxOutConnector[9] = fifoOut[24][9];
              muxOutConnector[10] = fifoOut[25][9];
              muxOutConnector[11] = fifoOut[0][8];
              muxOutConnector[12] = fifoOut[1][8];
              muxOutConnector[13] = fifoOut[2][8];
              muxOutConnector[14] = fifoOut[3][8];
              muxOutConnector[15] = fifoOut[4][8];
              muxOutConnector[16] = fifoOut[5][8];
              muxOutConnector[17] = fifoOut[6][8];
              muxOutConnector[18] = fifoOut[7][8];
              muxOutConnector[19] = fifoOut[8][8];
              muxOutConnector[20] = fifoOut[9][8];
              muxOutConnector[21] = fifoOut[10][8];
              muxOutConnector[22] = fifoOut[11][8];
              muxOutConnector[23] = fifoOut[12][8];
              muxOutConnector[24] = fifoOut[13][8];
              muxOutConnector[25] = fifoOut[14][8];
              muxOutConnector[26] = fifoOut[15][1];
              muxOutConnector[27] = fifoOut[16][1];
              muxOutConnector[28] = fifoOut[17][1];
              muxOutConnector[29] = fifoOut[18][1];
              muxOutConnector[30] = fifoOut[19][1];
              muxOutConnector[31] = fifoOut[20][1];
              muxOutConnector[32] = fifoOut[21][1];
              muxOutConnector[33] = fifoOut[22][1];
              muxOutConnector[34] = fifoOut[23][1];
              muxOutConnector[35] = fifoOut[24][1];
              muxOutConnector[36] = fifoOut[25][1];
              muxOutConnector[37] = fifoOut[0][0];
              muxOutConnector[38] = fifoOut[1][0];
              muxOutConnector[39] = fifoOut[2][0];
              muxOutConnector[40] = fifoOut[3][0];
              muxOutConnector[41] = fifoOut[4][0];
              muxOutConnector[42] = fifoOut[5][0];
              muxOutConnector[43] = fifoOut[6][0];
              muxOutConnector[44] = fifoOut[7][0];
              muxOutConnector[45] = fifoOut[8][0];
              muxOutConnector[46] = fifoOut[9][0];
              muxOutConnector[47] = fifoOut[10][0];
              muxOutConnector[48] = fifoOut[11][0];
              muxOutConnector[49] = fifoOut[12][0];
              muxOutConnector[50] = fifoOut[13][0];
              muxOutConnector[51] = fifoOut[14][0];
       end
       3: begin
              muxOutConnector[0] = fifoOut[15][9];
              muxOutConnector[1] = fifoOut[16][9];
              muxOutConnector[2] = fifoOut[17][9];
              muxOutConnector[3] = fifoOut[18][9];
              muxOutConnector[4] = fifoOut[19][9];
              muxOutConnector[5] = fifoOut[20][9];
              muxOutConnector[6] = fifoOut[21][9];
              muxOutConnector[7] = fifoOut[22][9];
              muxOutConnector[8] = fifoOut[23][9];
              muxOutConnector[9] = fifoOut[24][9];
              muxOutConnector[10] = fifoOut[25][9];
              muxOutConnector[11] = fifoOut[0][8];
              muxOutConnector[12] = fifoOut[1][8];
              muxOutConnector[13] = fifoOut[2][8];
              muxOutConnector[14] = fifoOut[3][8];
              muxOutConnector[15] = fifoOut[4][8];
              muxOutConnector[16] = fifoOut[5][8];
              muxOutConnector[17] = fifoOut[6][8];
              muxOutConnector[18] = fifoOut[7][8];
              muxOutConnector[19] = fifoOut[8][8];
              muxOutConnector[20] = fifoOut[9][8];
              muxOutConnector[21] = fifoOut[10][8];
              muxOutConnector[22] = fifoOut[11][8];
              muxOutConnector[23] = fifoOut[12][8];
              muxOutConnector[24] = fifoOut[13][8];
              muxOutConnector[25] = fifoOut[14][8];
              muxOutConnector[26] = fifoOut[15][1];
              muxOutConnector[27] = fifoOut[16][1];
              muxOutConnector[28] = fifoOut[17][1];
              muxOutConnector[29] = fifoOut[18][1];
              muxOutConnector[30] = fifoOut[19][1];
              muxOutConnector[31] = fifoOut[20][1];
              muxOutConnector[32] = fifoOut[21][1];
              muxOutConnector[33] = fifoOut[22][1];
              muxOutConnector[34] = fifoOut[23][1];
              muxOutConnector[35] = fifoOut[24][1];
              muxOutConnector[36] = fifoOut[25][1];
              muxOutConnector[37] = fifoOut[0][0];
              muxOutConnector[38] = fifoOut[1][0];
              muxOutConnector[39] = fifoOut[2][0];
              muxOutConnector[40] = fifoOut[3][0];
              muxOutConnector[41] = fifoOut[4][0];
              muxOutConnector[42] = fifoOut[5][0];
              muxOutConnector[43] = fifoOut[6][0];
              muxOutConnector[44] = fifoOut[7][0];
              muxOutConnector[45] = fifoOut[8][0];
              muxOutConnector[46] = fifoOut[9][0];
              muxOutConnector[47] = fifoOut[10][0];
              muxOutConnector[48] = fifoOut[11][0];
              muxOutConnector[49] = fifoOut[12][0];
              muxOutConnector[50] = fifoOut[13][0];
              muxOutConnector[51] = fifoOut[14][0];
       end
       4: begin
              muxOutConnector[0] = fifoOut[15][9];
              muxOutConnector[1] = fifoOut[16][9];
              muxOutConnector[2] = fifoOut[17][9];
              muxOutConnector[3] = fifoOut[18][9];
              muxOutConnector[4] = fifoOut[19][9];
              muxOutConnector[5] = fifoOut[20][9];
              muxOutConnector[6] = fifoOut[21][9];
              muxOutConnector[7] = fifoOut[22][9];
              muxOutConnector[8] = fifoOut[23][9];
              muxOutConnector[9] = fifoOut[24][9];
              muxOutConnector[10] = fifoOut[25][9];
              muxOutConnector[11] = fifoOut[0][8];
              muxOutConnector[12] = fifoOut[1][8];
              muxOutConnector[13] = fifoOut[2][8];
              muxOutConnector[14] = fifoOut[3][8];
              muxOutConnector[15] = fifoOut[4][8];
              muxOutConnector[16] = fifoOut[5][8];
              muxOutConnector[17] = fifoOut[6][8];
              muxOutConnector[18] = fifoOut[7][8];
              muxOutConnector[19] = fifoOut[8][8];
              muxOutConnector[20] = fifoOut[9][8];
              muxOutConnector[21] = fifoOut[10][8];
              muxOutConnector[22] = fifoOut[11][8];
              muxOutConnector[23] = fifoOut[12][8];
              muxOutConnector[24] = fifoOut[13][8];
              muxOutConnector[25] = fifoOut[14][8];
              muxOutConnector[26] = fifoOut[15][1];
              muxOutConnector[27] = fifoOut[16][1];
              muxOutConnector[28] = fifoOut[17][1];
              muxOutConnector[29] = fifoOut[18][1];
              muxOutConnector[30] = fifoOut[19][1];
              muxOutConnector[31] = fifoOut[20][1];
              muxOutConnector[32] = fifoOut[21][1];
              muxOutConnector[33] = fifoOut[22][1];
              muxOutConnector[34] = fifoOut[23][1];
              muxOutConnector[35] = fifoOut[24][1];
              muxOutConnector[36] = fifoOut[25][1];
              muxOutConnector[37] = fifoOut[0][0];
              muxOutConnector[38] = fifoOut[1][0];
              muxOutConnector[39] = fifoOut[2][0];
              muxOutConnector[40] = fifoOut[3][0];
              muxOutConnector[41] = fifoOut[4][0];
              muxOutConnector[42] = fifoOut[5][0];
              muxOutConnector[43] = fifoOut[6][0];
              muxOutConnector[44] = fifoOut[7][0];
              muxOutConnector[45] = fifoOut[8][0];
              muxOutConnector[46] = fifoOut[9][0];
              muxOutConnector[47] = fifoOut[10][0];
              muxOutConnector[48] = fifoOut[11][0];
              muxOutConnector[49] = fifoOut[12][0];
              muxOutConnector[50] = fifoOut[13][0];
              muxOutConnector[51] = fifoOut[14][0];
       end
       5: begin
              muxOutConnector[0] = fifoOut[15][9];
              muxOutConnector[1] = fifoOut[16][9];
              muxOutConnector[2] = fifoOut[17][9];
              muxOutConnector[3] = fifoOut[18][9];
              muxOutConnector[4] = fifoOut[19][9];
              muxOutConnector[5] = fifoOut[20][9];
              muxOutConnector[6] = fifoOut[21][9];
              muxOutConnector[7] = fifoOut[22][9];
              muxOutConnector[8] = fifoOut[23][9];
              muxOutConnector[9] = fifoOut[24][9];
              muxOutConnector[10] = fifoOut[25][9];
              muxOutConnector[11] = fifoOut[0][8];
              muxOutConnector[12] = fifoOut[1][8];
              muxOutConnector[13] = fifoOut[2][8];
              muxOutConnector[14] = fifoOut[3][8];
              muxOutConnector[15] = fifoOut[4][8];
              muxOutConnector[16] = fifoOut[5][8];
              muxOutConnector[17] = fifoOut[6][8];
              muxOutConnector[18] = fifoOut[7][8];
              muxOutConnector[19] = fifoOut[8][8];
              muxOutConnector[20] = fifoOut[9][8];
              muxOutConnector[21] = fifoOut[10][8];
              muxOutConnector[22] = fifoOut[11][8];
              muxOutConnector[23] = fifoOut[12][8];
              muxOutConnector[24] = fifoOut[13][8];
              muxOutConnector[25] = fifoOut[14][8];
              muxOutConnector[26] = fifoOut[15][1];
              muxOutConnector[27] = fifoOut[16][1];
              muxOutConnector[28] = fifoOut[17][1];
              muxOutConnector[29] = fifoOut[18][1];
              muxOutConnector[30] = fifoOut[19][1];
              muxOutConnector[31] = fifoOut[20][1];
              muxOutConnector[32] = fifoOut[21][1];
              muxOutConnector[33] = fifoOut[22][1];
              muxOutConnector[34] = fifoOut[23][1];
              muxOutConnector[35] = fifoOut[24][1];
              muxOutConnector[36] = fifoOut[25][1];
              muxOutConnector[37] = fifoOut[0][0];
              muxOutConnector[38] = fifoOut[1][0];
              muxOutConnector[39] = fifoOut[2][0];
              muxOutConnector[40] = fifoOut[3][0];
              muxOutConnector[41] = fifoOut[4][0];
              muxOutConnector[42] = fifoOut[5][0];
              muxOutConnector[43] = fifoOut[6][0];
              muxOutConnector[44] = fifoOut[7][0];
              muxOutConnector[45] = fifoOut[8][0];
              muxOutConnector[46] = fifoOut[9][0];
              muxOutConnector[47] = fifoOut[10][0];
              muxOutConnector[48] = fifoOut[11][0];
              muxOutConnector[49] = fifoOut[12][0];
              muxOutConnector[50] = fifoOut[13][0];
              muxOutConnector[51] = fifoOut[14][0];
       end
       6: begin
              muxOutConnector[0] = fifoOut[15][9];
              muxOutConnector[1] = fifoOut[16][9];
              muxOutConnector[2] = fifoOut[17][9];
              muxOutConnector[3] = fifoOut[18][9];
              muxOutConnector[4] = fifoOut[19][9];
              muxOutConnector[5] = fifoOut[20][9];
              muxOutConnector[6] = fifoOut[21][9];
              muxOutConnector[7] = fifoOut[22][9];
              muxOutConnector[8] = fifoOut[23][9];
              muxOutConnector[9] = fifoOut[24][9];
              muxOutConnector[10] = fifoOut[25][9];
              muxOutConnector[11] = fifoOut[0][8];
              muxOutConnector[12] = fifoOut[1][8];
              muxOutConnector[13] = fifoOut[2][8];
              muxOutConnector[14] = fifoOut[3][8];
              muxOutConnector[15] = fifoOut[4][8];
              muxOutConnector[16] = fifoOut[5][8];
              muxOutConnector[17] = fifoOut[6][8];
              muxOutConnector[18] = fifoOut[7][8];
              muxOutConnector[19] = fifoOut[8][8];
              muxOutConnector[20] = fifoOut[9][8];
              muxOutConnector[21] = fifoOut[10][8];
              muxOutConnector[22] = fifoOut[11][8];
              muxOutConnector[23] = fifoOut[12][8];
              muxOutConnector[24] = fifoOut[13][8];
              muxOutConnector[25] = fifoOut[14][8];
              muxOutConnector[26] = fifoOut[15][1];
              muxOutConnector[27] = fifoOut[16][1];
              muxOutConnector[28] = fifoOut[17][1];
              muxOutConnector[29] = fifoOut[18][1];
              muxOutConnector[30] = fifoOut[19][1];
              muxOutConnector[31] = fifoOut[20][1];
              muxOutConnector[32] = fifoOut[21][1];
              muxOutConnector[33] = fifoOut[22][1];
              muxOutConnector[34] = fifoOut[23][1];
              muxOutConnector[35] = fifoOut[24][1];
              muxOutConnector[36] = fifoOut[25][1];
              muxOutConnector[37] = fifoOut[0][0];
              muxOutConnector[38] = fifoOut[1][0];
              muxOutConnector[39] = fifoOut[2][0];
              muxOutConnector[40] = fifoOut[3][0];
              muxOutConnector[41] = fifoOut[4][0];
              muxOutConnector[42] = fifoOut[5][0];
              muxOutConnector[43] = fifoOut[6][0];
              muxOutConnector[44] = fifoOut[7][0];
              muxOutConnector[45] = fifoOut[8][0];
              muxOutConnector[46] = fifoOut[9][0];
              muxOutConnector[47] = fifoOut[10][0];
              muxOutConnector[48] = fifoOut[11][0];
              muxOutConnector[49] = fifoOut[12][0];
              muxOutConnector[50] = fifoOut[13][0];
              muxOutConnector[51] = fifoOut[14][0];
       end
       7: begin
              muxOutConnector[0] = fifoOut[15][9];
              muxOutConnector[1] = fifoOut[16][9];
              muxOutConnector[2] = fifoOut[17][9];
              muxOutConnector[3] = fifoOut[18][9];
              muxOutConnector[4] = fifoOut[19][9];
              muxOutConnector[5] = fifoOut[20][9];
              muxOutConnector[6] = fifoOut[21][9];
              muxOutConnector[7] = fifoOut[22][9];
              muxOutConnector[8] = fifoOut[23][9];
              muxOutConnector[9] = fifoOut[24][9];
              muxOutConnector[10] = fifoOut[25][9];
              muxOutConnector[11] = fifoOut[0][8];
              muxOutConnector[12] = fifoOut[1][8];
              muxOutConnector[13] = fifoOut[2][8];
              muxOutConnector[14] = fifoOut[3][8];
              muxOutConnector[15] = fifoOut[4][8];
              muxOutConnector[16] = fifoOut[5][8];
              muxOutConnector[17] = fifoOut[6][8];
              muxOutConnector[18] = fifoOut[7][8];
              muxOutConnector[19] = fifoOut[8][8];
              muxOutConnector[20] = fifoOut[9][8];
              muxOutConnector[21] = fifoOut[10][8];
              muxOutConnector[22] = fifoOut[11][8];
              muxOutConnector[23] = fifoOut[12][8];
              muxOutConnector[24] = fifoOut[13][8];
              muxOutConnector[25] = fifoOut[14][8];
              muxOutConnector[26] = fifoOut[15][1];
              muxOutConnector[27] = fifoOut[16][1];
              muxOutConnector[28] = fifoOut[17][1];
              muxOutConnector[29] = fifoOut[18][1];
              muxOutConnector[30] = fifoOut[19][1];
              muxOutConnector[31] = fifoOut[20][1];
              muxOutConnector[32] = fifoOut[21][1];
              muxOutConnector[33] = fifoOut[22][1];
              muxOutConnector[34] = fifoOut[23][1];
              muxOutConnector[35] = fifoOut[24][1];
              muxOutConnector[36] = fifoOut[25][1];
              muxOutConnector[37] = fifoOut[0][0];
              muxOutConnector[38] = fifoOut[1][0];
              muxOutConnector[39] = fifoOut[2][0];
              muxOutConnector[40] = fifoOut[3][0];
              muxOutConnector[41] = fifoOut[4][0];
              muxOutConnector[42] = fifoOut[5][0];
              muxOutConnector[43] = fifoOut[6][0];
              muxOutConnector[44] = fifoOut[7][0];
              muxOutConnector[45] = fifoOut[8][0];
              muxOutConnector[46] = fifoOut[9][0];
              muxOutConnector[47] = fifoOut[10][0];
              muxOutConnector[48] = fifoOut[11][0];
              muxOutConnector[49] = fifoOut[12][0];
              muxOutConnector[50] = fifoOut[13][0];
              muxOutConnector[51] = fifoOut[14][0];
       end
       8: begin
              muxOutConnector[0] = fifoOut[15][9];
              muxOutConnector[1] = fifoOut[16][9];
              muxOutConnector[2] = fifoOut[17][9];
              muxOutConnector[3] = fifoOut[18][9];
              muxOutConnector[4] = fifoOut[19][9];
              muxOutConnector[5] = fifoOut[20][9];
              muxOutConnector[6] = fifoOut[21][9];
              muxOutConnector[7] = fifoOut[22][9];
              muxOutConnector[8] = fifoOut[23][9];
              muxOutConnector[9] = fifoOut[24][9];
              muxOutConnector[10] = fifoOut[25][9];
              muxOutConnector[11] = fifoOut[0][8];
              muxOutConnector[12] = fifoOut[1][8];
              muxOutConnector[13] = fifoOut[2][8];
              muxOutConnector[14] = fifoOut[3][8];
              muxOutConnector[15] = fifoOut[4][8];
              muxOutConnector[16] = fifoOut[5][8];
              muxOutConnector[17] = fifoOut[6][8];
              muxOutConnector[18] = fifoOut[7][8];
              muxOutConnector[19] = fifoOut[8][8];
              muxOutConnector[20] = fifoOut[9][8];
              muxOutConnector[21] = fifoOut[10][8];
              muxOutConnector[22] = fifoOut[11][8];
              muxOutConnector[23] = fifoOut[12][8];
              muxOutConnector[24] = fifoOut[13][8];
              muxOutConnector[25] = fifoOut[14][8];
              muxOutConnector[26] = fifoOut[15][1];
              muxOutConnector[27] = fifoOut[16][1];
              muxOutConnector[28] = fifoOut[17][1];
              muxOutConnector[29] = fifoOut[18][1];
              muxOutConnector[30] = fifoOut[19][1];
              muxOutConnector[31] = fifoOut[20][1];
              muxOutConnector[32] = fifoOut[21][1];
              muxOutConnector[33] = fifoOut[22][1];
              muxOutConnector[34] = fifoOut[23][1];
              muxOutConnector[35] = fifoOut[24][1];
              muxOutConnector[36] = fifoOut[25][1];
              muxOutConnector[37] = fifoOut[0][0];
              muxOutConnector[38] = fifoOut[1][0];
              muxOutConnector[39] = fifoOut[2][0];
              muxOutConnector[40] = fifoOut[3][0];
              muxOutConnector[41] = fifoOut[4][0];
              muxOutConnector[42] = fifoOut[5][0];
              muxOutConnector[43] = fifoOut[6][0];
              muxOutConnector[44] = fifoOut[7][0];
              muxOutConnector[45] = fifoOut[8][0];
              muxOutConnector[46] = fifoOut[9][0];
              muxOutConnector[47] = fifoOut[10][0];
              muxOutConnector[48] = fifoOut[11][0];
              muxOutConnector[49] = fifoOut[12][0];
              muxOutConnector[50] = fifoOut[13][0];
              muxOutConnector[51] = fifoOut[14][0];
       end
       9: begin
              muxOutConnector[0] = fifoOut[15][9];
              muxOutConnector[1] = fifoOut[16][9];
              muxOutConnector[2] = fifoOut[33][5];
              muxOutConnector[3] = fifoOut[34][5];
              muxOutConnector[4] = fifoOut[35][5];
              muxOutConnector[5] = fifoOut[36][5];
              muxOutConnector[6] = fifoOut[37][5];
              muxOutConnector[7] = fifoOut[38][5];
              muxOutConnector[8] = fifoOut[39][5];
              muxOutConnector[9] = fifoOut[40][5];
              muxOutConnector[10] = fifoOut[41][5];
              muxOutConnector[11] = fifoOut[42][5];
              muxOutConnector[12] = fifoOut[43][5];
              muxOutConnector[13] = fifoOut[44][5];
              muxOutConnector[14] = fifoOut[45][5];
              muxOutConnector[15] = fifoOut[46][5];
              muxOutConnector[16] = fifoOut[47][5];
              muxOutConnector[17] = fifoOut[48][5];
              muxOutConnector[18] = fifoOut[49][5];
              muxOutConnector[19] = fifoOut[50][5];
              muxOutConnector[20] = fifoOut[51][5];
              muxOutConnector[21] = fifoOut[26][4];
              muxOutConnector[22] = fifoOut[27][4];
              muxOutConnector[23] = fifoOut[28][4];
              muxOutConnector[24] = fifoOut[29][4];
              muxOutConnector[25] = fifoOut[30][4];
              muxOutConnector[26] = fifoOut[15][1];
              muxOutConnector[27] = fifoOut[16][1];
              muxOutConnector[28] = fifoOut[17][1];
              muxOutConnector[29] = fifoOut[18][1];
              muxOutConnector[30] = fifoOut[19][1];
              muxOutConnector[31] = fifoOut[20][1];
              muxOutConnector[32] = fifoOut[21][1];
              muxOutConnector[33] = fifoOut[22][1];
              muxOutConnector[34] = fifoOut[23][1];
              muxOutConnector[35] = fifoOut[24][1];
              muxOutConnector[36] = fifoOut[25][1];
              muxOutConnector[37] = fifoOut[0][0];
              muxOutConnector[38] = fifoOut[1][0];
              muxOutConnector[39] = fifoOut[2][0];
              muxOutConnector[40] = fifoOut[3][0];
              muxOutConnector[41] = fifoOut[4][0];
              muxOutConnector[42] = fifoOut[5][0];
              muxOutConnector[43] = fifoOut[6][0];
              muxOutConnector[44] = fifoOut[7][0];
              muxOutConnector[45] = fifoOut[8][0];
              muxOutConnector[46] = fifoOut[9][0];
              muxOutConnector[47] = fifoOut[26][8];
              muxOutConnector[48] = fifoOut[27][8];
              muxOutConnector[49] = fifoOut[28][8];
              muxOutConnector[50] = fifoOut[29][8];
              muxOutConnector[51] = fifoOut[30][8];
       end
       10: begin
              muxOutConnector[0] = fifoOut[31][5];
              muxOutConnector[1] = fifoOut[32][5];
              muxOutConnector[2] = fifoOut[33][5];
              muxOutConnector[3] = fifoOut[34][5];
              muxOutConnector[4] = fifoOut[35][5];
              muxOutConnector[5] = fifoOut[36][5];
              muxOutConnector[6] = fifoOut[37][5];
              muxOutConnector[7] = fifoOut[38][5];
              muxOutConnector[8] = fifoOut[39][5];
              muxOutConnector[9] = fifoOut[40][5];
              muxOutConnector[10] = fifoOut[41][5];
              muxOutConnector[11] = fifoOut[42][5];
              muxOutConnector[12] = fifoOut[43][5];
              muxOutConnector[13] = fifoOut[44][5];
              muxOutConnector[14] = fifoOut[45][5];
              muxOutConnector[15] = fifoOut[46][5];
              muxOutConnector[16] = fifoOut[47][5];
              muxOutConnector[17] = fifoOut[48][5];
              muxOutConnector[18] = fifoOut[49][5];
              muxOutConnector[19] = fifoOut[50][5];
              muxOutConnector[20] = fifoOut[51][5];
              muxOutConnector[21] = fifoOut[26][4];
              muxOutConnector[22] = fifoOut[27][4];
              muxOutConnector[23] = fifoOut[28][4];
              muxOutConnector[24] = fifoOut[29][4];
              muxOutConnector[25] = fifoOut[30][4];
              muxOutConnector[26] = fifoOut[31][9];
              muxOutConnector[27] = fifoOut[32][9];
              muxOutConnector[28] = fifoOut[33][9];
              muxOutConnector[29] = fifoOut[34][9];
              muxOutConnector[30] = fifoOut[35][9];
              muxOutConnector[31] = fifoOut[36][9];
              muxOutConnector[32] = fifoOut[37][9];
              muxOutConnector[33] = fifoOut[38][9];
              muxOutConnector[34] = fifoOut[39][9];
              muxOutConnector[35] = fifoOut[40][9];
              muxOutConnector[36] = fifoOut[41][9];
              muxOutConnector[37] = fifoOut[42][9];
              muxOutConnector[38] = fifoOut[43][9];
              muxOutConnector[39] = fifoOut[44][9];
              muxOutConnector[40] = fifoOut[45][9];
              muxOutConnector[41] = fifoOut[46][9];
              muxOutConnector[42] = fifoOut[47][9];
              muxOutConnector[43] = fifoOut[48][9];
              muxOutConnector[44] = fifoOut[49][9];
              muxOutConnector[45] = fifoOut[50][9];
              muxOutConnector[46] = fifoOut[51][9];
              muxOutConnector[47] = fifoOut[26][8];
              muxOutConnector[48] = fifoOut[27][8];
              muxOutConnector[49] = fifoOut[28][8];
              muxOutConnector[50] = fifoOut[29][8];
              muxOutConnector[51] = fifoOut[30][8];
       end
       11: begin
              muxOutConnector[0] = fifoOut[31][5];
              muxOutConnector[1] = fifoOut[32][5];
              muxOutConnector[2] = fifoOut[33][5];
              muxOutConnector[3] = fifoOut[34][5];
              muxOutConnector[4] = fifoOut[35][5];
              muxOutConnector[5] = fifoOut[36][5];
              muxOutConnector[6] = fifoOut[37][5];
              muxOutConnector[7] = fifoOut[38][5];
              muxOutConnector[8] = fifoOut[39][5];
              muxOutConnector[9] = fifoOut[40][5];
              muxOutConnector[10] = fifoOut[41][5];
              muxOutConnector[11] = fifoOut[42][5];
              muxOutConnector[12] = fifoOut[43][5];
              muxOutConnector[13] = fifoOut[44][5];
              muxOutConnector[14] = fifoOut[45][5];
              muxOutConnector[15] = fifoOut[46][5];
              muxOutConnector[16] = fifoOut[47][5];
              muxOutConnector[17] = fifoOut[48][5];
              muxOutConnector[18] = fifoOut[49][5];
              muxOutConnector[19] = fifoOut[50][5];
              muxOutConnector[20] = fifoOut[51][5];
              muxOutConnector[21] = fifoOut[26][4];
              muxOutConnector[22] = fifoOut[27][4];
              muxOutConnector[23] = fifoOut[28][4];
              muxOutConnector[24] = fifoOut[29][4];
              muxOutConnector[25] = fifoOut[30][4];
              muxOutConnector[26] = fifoOut[31][9];
              muxOutConnector[27] = fifoOut[32][9];
              muxOutConnector[28] = fifoOut[33][9];
              muxOutConnector[29] = fifoOut[34][9];
              muxOutConnector[30] = fifoOut[35][9];
              muxOutConnector[31] = fifoOut[36][9];
              muxOutConnector[32] = fifoOut[37][9];
              muxOutConnector[33] = fifoOut[38][9];
              muxOutConnector[34] = fifoOut[39][9];
              muxOutConnector[35] = fifoOut[40][9];
              muxOutConnector[36] = fifoOut[41][9];
              muxOutConnector[37] = fifoOut[42][9];
              muxOutConnector[38] = fifoOut[43][9];
              muxOutConnector[39] = fifoOut[44][9];
              muxOutConnector[40] = fifoOut[45][9];
              muxOutConnector[41] = fifoOut[46][9];
              muxOutConnector[42] = fifoOut[47][9];
              muxOutConnector[43] = fifoOut[48][9];
              muxOutConnector[44] = fifoOut[49][9];
              muxOutConnector[45] = fifoOut[50][9];
              muxOutConnector[46] = fifoOut[51][9];
              muxOutConnector[47] = fifoOut[26][8];
              muxOutConnector[48] = fifoOut[27][8];
              muxOutConnector[49] = fifoOut[28][8];
              muxOutConnector[50] = fifoOut[29][8];
              muxOutConnector[51] = fifoOut[30][8];
       end
       12: begin
              muxOutConnector[0] = fifoOut[31][5];
              muxOutConnector[1] = fifoOut[32][5];
              muxOutConnector[2] = fifoOut[33][5];
              muxOutConnector[3] = fifoOut[34][5];
              muxOutConnector[4] = fifoOut[35][5];
              muxOutConnector[5] = fifoOut[36][5];
              muxOutConnector[6] = fifoOut[37][5];
              muxOutConnector[7] = fifoOut[38][5];
              muxOutConnector[8] = fifoOut[39][5];
              muxOutConnector[9] = fifoOut[40][5];
              muxOutConnector[10] = fifoOut[41][5];
              muxOutConnector[11] = fifoOut[42][5];
              muxOutConnector[12] = fifoOut[43][5];
              muxOutConnector[13] = fifoOut[44][5];
              muxOutConnector[14] = fifoOut[45][5];
              muxOutConnector[15] = fifoOut[46][5];
              muxOutConnector[16] = fifoOut[47][5];
              muxOutConnector[17] = fifoOut[48][5];
              muxOutConnector[18] = fifoOut[49][5];
              muxOutConnector[19] = fifoOut[50][5];
              muxOutConnector[20] = fifoOut[51][5];
              muxOutConnector[21] = fifoOut[26][4];
              muxOutConnector[22] = fifoOut[27][4];
              muxOutConnector[23] = fifoOut[28][4];
              muxOutConnector[24] = fifoOut[29][4];
              muxOutConnector[25] = fifoOut[30][4];
              muxOutConnector[26] = fifoOut[31][9];
              muxOutConnector[27] = fifoOut[32][9];
              muxOutConnector[28] = fifoOut[33][9];
              muxOutConnector[29] = fifoOut[34][9];
              muxOutConnector[30] = fifoOut[35][9];
              muxOutConnector[31] = fifoOut[36][9];
              muxOutConnector[32] = fifoOut[37][9];
              muxOutConnector[33] = fifoOut[38][9];
              muxOutConnector[34] = fifoOut[39][9];
              muxOutConnector[35] = fifoOut[40][9];
              muxOutConnector[36] = fifoOut[41][9];
              muxOutConnector[37] = fifoOut[42][9];
              muxOutConnector[38] = fifoOut[43][9];
              muxOutConnector[39] = fifoOut[44][9];
              muxOutConnector[40] = fifoOut[45][9];
              muxOutConnector[41] = fifoOut[46][9];
              muxOutConnector[42] = fifoOut[47][9];
              muxOutConnector[43] = fifoOut[48][9];
              muxOutConnector[44] = fifoOut[49][9];
              muxOutConnector[45] = fifoOut[50][9];
              muxOutConnector[46] = fifoOut[51][9];
              muxOutConnector[47] = fifoOut[26][8];
              muxOutConnector[48] = fifoOut[27][8];
              muxOutConnector[49] = fifoOut[28][8];
              muxOutConnector[50] = fifoOut[29][8];
              muxOutConnector[51] = fifoOut[30][8];
       end
       13: begin
              muxOutConnector[0] = fifoOut[31][5];
              muxOutConnector[1] = fifoOut[32][5];
              muxOutConnector[2] = fifoOut[33][5];
              muxOutConnector[3] = fifoOut[34][5];
              muxOutConnector[4] = fifoOut[35][5];
              muxOutConnector[5] = fifoOut[36][5];
              muxOutConnector[6] = fifoOut[37][5];
              muxOutConnector[7] = fifoOut[38][5];
              muxOutConnector[8] = fifoOut[39][5];
              muxOutConnector[9] = fifoOut[40][5];
              muxOutConnector[10] = fifoOut[41][5];
              muxOutConnector[11] = fifoOut[42][5];
              muxOutConnector[12] = fifoOut[43][5];
              muxOutConnector[13] = fifoOut[44][5];
              muxOutConnector[14] = fifoOut[45][5];
              muxOutConnector[15] = fifoOut[46][5];
              muxOutConnector[16] = fifoOut[47][5];
              muxOutConnector[17] = fifoOut[48][5];
              muxOutConnector[18] = fifoOut[49][5];
              muxOutConnector[19] = fifoOut[50][5];
              muxOutConnector[20] = fifoOut[51][5];
              muxOutConnector[21] = fifoOut[26][4];
              muxOutConnector[22] = fifoOut[27][4];
              muxOutConnector[23] = fifoOut[28][4];
              muxOutConnector[24] = fifoOut[29][4];
              muxOutConnector[25] = fifoOut[30][4];
              muxOutConnector[26] = fifoOut[31][9];
              muxOutConnector[27] = fifoOut[32][9];
              muxOutConnector[28] = fifoOut[33][9];
              muxOutConnector[29] = fifoOut[34][9];
              muxOutConnector[30] = fifoOut[35][9];
              muxOutConnector[31] = fifoOut[36][9];
              muxOutConnector[32] = fifoOut[37][9];
              muxOutConnector[33] = fifoOut[38][9];
              muxOutConnector[34] = fifoOut[39][9];
              muxOutConnector[35] = fifoOut[40][9];
              muxOutConnector[36] = fifoOut[41][9];
              muxOutConnector[37] = fifoOut[42][9];
              muxOutConnector[38] = fifoOut[43][9];
              muxOutConnector[39] = fifoOut[44][9];
              muxOutConnector[40] = fifoOut[45][9];
              muxOutConnector[41] = fifoOut[46][9];
              muxOutConnector[42] = fifoOut[47][9];
              muxOutConnector[43] = fifoOut[48][9];
              muxOutConnector[44] = fifoOut[49][9];
              muxOutConnector[45] = fifoOut[50][9];
              muxOutConnector[46] = fifoOut[51][9];
              muxOutConnector[47] = fifoOut[26][8];
              muxOutConnector[48] = fifoOut[27][8];
              muxOutConnector[49] = fifoOut[28][8];
              muxOutConnector[50] = fifoOut[29][8];
              muxOutConnector[51] = fifoOut[30][8];
       end
       14: begin
              muxOutConnector[0] = fifoOut[31][5];
              muxOutConnector[1] = fifoOut[32][5];
              muxOutConnector[2] = fifoOut[33][5];
              muxOutConnector[3] = fifoOut[34][5];
              muxOutConnector[4] = fifoOut[35][5];
              muxOutConnector[5] = fifoOut[36][5];
              muxOutConnector[6] = fifoOut[37][5];
              muxOutConnector[7] = fifoOut[38][5];
              muxOutConnector[8] = fifoOut[39][5];
              muxOutConnector[9] = fifoOut[40][5];
              muxOutConnector[10] = fifoOut[41][5];
              muxOutConnector[11] = fifoOut[42][5];
              muxOutConnector[12] = fifoOut[43][5];
              muxOutConnector[13] = fifoOut[44][5];
              muxOutConnector[14] = fifoOut[45][5];
              muxOutConnector[15] = fifoOut[46][5];
              muxOutConnector[16] = fifoOut[47][5];
              muxOutConnector[17] = fifoOut[48][5];
              muxOutConnector[18] = fifoOut[49][5];
              muxOutConnector[19] = fifoOut[50][5];
              muxOutConnector[20] = fifoOut[51][5];
              muxOutConnector[21] = fifoOut[26][4];
              muxOutConnector[22] = fifoOut[27][4];
              muxOutConnector[23] = fifoOut[28][4];
              muxOutConnector[24] = fifoOut[29][4];
              muxOutConnector[25] = fifoOut[30][4];
              muxOutConnector[26] = fifoOut[31][9];
              muxOutConnector[27] = fifoOut[32][9];
              muxOutConnector[28] = fifoOut[33][9];
              muxOutConnector[29] = fifoOut[34][9];
              muxOutConnector[30] = fifoOut[35][9];
              muxOutConnector[31] = fifoOut[36][9];
              muxOutConnector[32] = fifoOut[37][9];
              muxOutConnector[33] = fifoOut[38][9];
              muxOutConnector[34] = fifoOut[39][9];
              muxOutConnector[35] = fifoOut[40][9];
              muxOutConnector[36] = fifoOut[41][9];
              muxOutConnector[37] = fifoOut[42][9];
              muxOutConnector[38] = fifoOut[43][9];
              muxOutConnector[39] = fifoOut[44][9];
              muxOutConnector[40] = fifoOut[45][9];
              muxOutConnector[41] = fifoOut[46][9];
              muxOutConnector[42] = fifoOut[47][9];
              muxOutConnector[43] = fifoOut[48][9];
              muxOutConnector[44] = fifoOut[49][9];
              muxOutConnector[45] = fifoOut[50][9];
              muxOutConnector[46] = fifoOut[51][9];
              muxOutConnector[47] = fifoOut[26][8];
              muxOutConnector[48] = fifoOut[27][8];
              muxOutConnector[49] = fifoOut[28][8];
              muxOutConnector[50] = fifoOut[29][8];
              muxOutConnector[51] = fifoOut[30][8];
       end
       15: begin
              muxOutConnector[0] = fifoOut[31][5];
              muxOutConnector[1] = fifoOut[32][5];
              muxOutConnector[2] = fifoOut[33][5];
              muxOutConnector[3] = fifoOut[34][5];
              muxOutConnector[4] = fifoOut[35][5];
              muxOutConnector[5] = fifoOut[36][5];
              muxOutConnector[6] = fifoOut[37][5];
              muxOutConnector[7] = fifoOut[38][5];
              muxOutConnector[8] = fifoOut[39][5];
              muxOutConnector[9] = fifoOut[40][5];
              muxOutConnector[10] = fifoOut[41][5];
              muxOutConnector[11] = fifoOut[42][5];
              muxOutConnector[12] = fifoOut[43][5];
              muxOutConnector[13] = fifoOut[44][5];
              muxOutConnector[14] = fifoOut[45][5];
              muxOutConnector[15] = fifoOut[46][5];
              muxOutConnector[16] = fifoOut[47][5];
              muxOutConnector[17] = fifoOut[48][5];
              muxOutConnector[18] = fifoOut[49][5];
              muxOutConnector[19] = fifoOut[50][5];
              muxOutConnector[20] = fifoOut[51][5];
              muxOutConnector[21] = fifoOut[26][4];
              muxOutConnector[22] = fifoOut[27][4];
              muxOutConnector[23] = fifoOut[28][4];
              muxOutConnector[24] = fifoOut[29][4];
              muxOutConnector[25] = fifoOut[30][4];
              muxOutConnector[26] = fifoOut[31][9];
              muxOutConnector[27] = fifoOut[32][9];
              muxOutConnector[28] = fifoOut[33][9];
              muxOutConnector[29] = fifoOut[34][9];
              muxOutConnector[30] = fifoOut[35][9];
              muxOutConnector[31] = fifoOut[36][9];
              muxOutConnector[32] = fifoOut[37][9];
              muxOutConnector[33] = fifoOut[38][9];
              muxOutConnector[34] = fifoOut[39][9];
              muxOutConnector[35] = fifoOut[40][9];
              muxOutConnector[36] = fifoOut[41][9];
              muxOutConnector[37] = fifoOut[42][9];
              muxOutConnector[38] = fifoOut[43][9];
              muxOutConnector[39] = fifoOut[44][9];
              muxOutConnector[40] = fifoOut[45][9];
              muxOutConnector[41] = fifoOut[46][9];
              muxOutConnector[42] = fifoOut[47][9];
              muxOutConnector[43] = fifoOut[48][9];
              muxOutConnector[44] = fifoOut[49][9];
              muxOutConnector[45] = fifoOut[50][9];
              muxOutConnector[46] = fifoOut[51][9];
              muxOutConnector[47] = fifoOut[26][8];
              muxOutConnector[48] = fifoOut[27][8];
              muxOutConnector[49] = fifoOut[28][8];
              muxOutConnector[50] = fifoOut[29][8];
              muxOutConnector[51] = fifoOut[30][8];
       end
       16: begin
              muxOutConnector[0] = fifoOut[31][5];
              muxOutConnector[1] = fifoOut[32][5];
              muxOutConnector[2] = fifoOut[33][5];
              muxOutConnector[3] = fifoOut[34][5];
              muxOutConnector[4] = fifoOut[35][5];
              muxOutConnector[5] = fifoOut[36][5];
              muxOutConnector[6] = fifoOut[37][5];
              muxOutConnector[7] = fifoOut[38][5];
              muxOutConnector[8] = fifoOut[39][5];
              muxOutConnector[9] = fifoOut[40][5];
              muxOutConnector[10] = fifoOut[41][5];
              muxOutConnector[11] = fifoOut[42][5];
              muxOutConnector[12] = fifoOut[43][5];
              muxOutConnector[13] = fifoOut[44][5];
              muxOutConnector[14] = fifoOut[45][5];
              muxOutConnector[15] = fifoOut[46][5];
              muxOutConnector[16] = fifoOut[47][5];
              muxOutConnector[17] = fifoOut[48][5];
              muxOutConnector[18] = fifoOut[49][5];
              muxOutConnector[19] = fifoOut[50][5];
              muxOutConnector[20] = fifoOut[51][5];
              muxOutConnector[21] = fifoOut[26][4];
              muxOutConnector[22] = fifoOut[27][4];
              muxOutConnector[23] = fifoOut[28][4];
              muxOutConnector[24] = fifoOut[29][4];
              muxOutConnector[25] = fifoOut[30][4];
              muxOutConnector[26] = fifoOut[31][9];
              muxOutConnector[27] = fifoOut[32][9];
              muxOutConnector[28] = fifoOut[33][9];
              muxOutConnector[29] = fifoOut[34][9];
              muxOutConnector[30] = fifoOut[35][9];
              muxOutConnector[31] = fifoOut[36][9];
              muxOutConnector[32] = fifoOut[37][9];
              muxOutConnector[33] = fifoOut[38][9];
              muxOutConnector[34] = fifoOut[39][9];
              muxOutConnector[35] = fifoOut[40][9];
              muxOutConnector[36] = fifoOut[41][9];
              muxOutConnector[37] = fifoOut[42][9];
              muxOutConnector[38] = fifoOut[43][9];
              muxOutConnector[39] = fifoOut[44][9];
              muxOutConnector[40] = fifoOut[45][9];
              muxOutConnector[41] = fifoOut[46][9];
              muxOutConnector[42] = fifoOut[47][9];
              muxOutConnector[43] = fifoOut[48][9];
              muxOutConnector[44] = fifoOut[49][9];
              muxOutConnector[45] = fifoOut[50][9];
              muxOutConnector[46] = fifoOut[51][9];
              muxOutConnector[47] = fifoOut[26][8];
              muxOutConnector[48] = fifoOut[27][8];
              muxOutConnector[49] = fifoOut[28][8];
              muxOutConnector[50] = fifoOut[29][8];
              muxOutConnector[51] = fifoOut[30][8];
       end
       17: begin
              muxOutConnector[0] = fifoOut[31][5];
              muxOutConnector[1] = fifoOut[32][5];
              muxOutConnector[2] = fifoOut[33][5];
              muxOutConnector[3] = fifoOut[34][5];
              muxOutConnector[4] = fifoOut[35][5];
              muxOutConnector[5] = fifoOut[36][5];
              muxOutConnector[6] = fifoOut[37][5];
              muxOutConnector[7] = fifoOut[38][5];
              muxOutConnector[8] = fifoOut[39][5];
              muxOutConnector[9] = fifoOut[40][5];
              muxOutConnector[10] = fifoOut[41][5];
              muxOutConnector[11] = fifoOut[42][5];
              muxOutConnector[12] = fifoOut[10][4];
              muxOutConnector[13] = fifoOut[11][4];
              muxOutConnector[14] = fifoOut[12][4];
              muxOutConnector[15] = fifoOut[13][4];
              muxOutConnector[16] = fifoOut[14][4];
              muxOutConnector[17] = fifoOut[15][4];
              muxOutConnector[18] = fifoOut[16][4];
              muxOutConnector[19] = fifoOut[17][4];
              muxOutConnector[20] = fifoOut[18][4];
              muxOutConnector[21] = fifoOut[19][4];
              muxOutConnector[22] = fifoOut[20][4];
              muxOutConnector[23] = fifoOut[21][4];
              muxOutConnector[24] = fifoOut[22][4];
              muxOutConnector[25] = fifoOut[23][4];
              muxOutConnector[26] = fifoOut[31][9];
              muxOutConnector[27] = fifoOut[32][9];
              muxOutConnector[28] = fifoOut[33][9];
              muxOutConnector[29] = fifoOut[34][9];
              muxOutConnector[30] = fifoOut[35][9];
              muxOutConnector[31] = fifoOut[36][9];
              muxOutConnector[32] = fifoOut[37][9];
              muxOutConnector[33] = fifoOut[38][9];
              muxOutConnector[34] = fifoOut[39][9];
              muxOutConnector[35] = fifoOut[40][9];
              muxOutConnector[36] = fifoOut[41][9];
              muxOutConnector[37] = fifoOut[42][9];
              muxOutConnector[38] = fifoOut[43][9];
              muxOutConnector[39] = fifoOut[44][9];
              muxOutConnector[40] = fifoOut[45][9];
              muxOutConnector[41] = fifoOut[46][9];
              muxOutConnector[42] = fifoOut[47][9];
              muxOutConnector[43] = fifoOut[48][9];
              muxOutConnector[44] = fifoOut[49][9];
              muxOutConnector[45] = fifoOut[50][9];
              muxOutConnector[46] = fifoOut[51][9];
              muxOutConnector[47] = fifoOut[26][8];
              muxOutConnector[48] = fifoOut[27][8];
              muxOutConnector[49] = fifoOut[28][8];
              muxOutConnector[50] = fifoOut[29][8];
              muxOutConnector[51] = fifoOut[30][8];
       end
       18: begin
              muxOutConnector[0] = fifoOut[24][5];
              muxOutConnector[1] = fifoOut[25][5];
              muxOutConnector[2] = fifoOut[0][4];
              muxOutConnector[3] = fifoOut[1][4];
              muxOutConnector[4] = fifoOut[2][4];
              muxOutConnector[5] = fifoOut[3][4];
              muxOutConnector[6] = fifoOut[4][4];
              muxOutConnector[7] = fifoOut[5][4];
              muxOutConnector[8] = fifoOut[6][4];
              muxOutConnector[9] = fifoOut[7][4];
              muxOutConnector[10] = fifoOut[8][4];
              muxOutConnector[11] = fifoOut[9][4];
              muxOutConnector[12] = fifoOut[10][4];
              muxOutConnector[13] = fifoOut[11][4];
              muxOutConnector[14] = fifoOut[12][4];
              muxOutConnector[15] = fifoOut[13][4];
              muxOutConnector[16] = fifoOut[14][4];
              muxOutConnector[17] = fifoOut[15][4];
              muxOutConnector[18] = fifoOut[16][4];
              muxOutConnector[19] = fifoOut[17][4];
              muxOutConnector[20] = fifoOut[18][4];
              muxOutConnector[21] = fifoOut[19][4];
              muxOutConnector[22] = fifoOut[20][4];
              muxOutConnector[23] = fifoOut[21][4];
              muxOutConnector[24] = fifoOut[22][4];
              muxOutConnector[25] = fifoOut[23][4];
              muxOutConnector[26] = fifoOut[31][9];
              muxOutConnector[27] = fifoOut[32][9];
              muxOutConnector[28] = fifoOut[33][9];
              muxOutConnector[29] = fifoOut[34][9];
              muxOutConnector[30] = fifoOut[35][9];
              muxOutConnector[31] = fifoOut[36][9];
              muxOutConnector[32] = fifoOut[37][9];
              muxOutConnector[33] = fifoOut[38][9];
              muxOutConnector[34] = fifoOut[39][9];
              muxOutConnector[35] = fifoOut[40][9];
              muxOutConnector[36] = fifoOut[41][9];
              muxOutConnector[37] = fifoOut[42][9];
              muxOutConnector[38] = fifoOut[43][9];
              muxOutConnector[39] = fifoOut[44][9];
              muxOutConnector[40] = fifoOut[45][9];
              muxOutConnector[41] = fifoOut[46][9];
              muxOutConnector[42] = fifoOut[47][9];
              muxOutConnector[43] = fifoOut[48][9];
              muxOutConnector[44] = fifoOut[49][9];
              muxOutConnector[45] = fifoOut[50][9];
              muxOutConnector[46] = fifoOut[51][9];
              muxOutConnector[47] = fifoOut[26][8];
              muxOutConnector[48] = fifoOut[27][8];
              muxOutConnector[49] = fifoOut[28][8];
              muxOutConnector[50] = fifoOut[29][8];
              muxOutConnector[51] = fifoOut[30][8];
       end
       19: begin
              muxOutConnector[0] = fifoOut[24][5];
              muxOutConnector[1] = fifoOut[25][5];
              muxOutConnector[2] = fifoOut[0][4];
              muxOutConnector[3] = fifoOut[1][4];
              muxOutConnector[4] = fifoOut[2][4];
              muxOutConnector[5] = fifoOut[3][4];
              muxOutConnector[6] = fifoOut[4][4];
              muxOutConnector[7] = fifoOut[5][4];
              muxOutConnector[8] = fifoOut[6][4];
              muxOutConnector[9] = fifoOut[7][4];
              muxOutConnector[10] = fifoOut[8][4];
              muxOutConnector[11] = fifoOut[9][4];
              muxOutConnector[12] = fifoOut[10][4];
              muxOutConnector[13] = fifoOut[11][4];
              muxOutConnector[14] = fifoOut[12][4];
              muxOutConnector[15] = fifoOut[13][4];
              muxOutConnector[16] = fifoOut[14][4];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[31][9];
              muxOutConnector[27] = fifoOut[32][9];
              muxOutConnector[28] = fifoOut[33][9];
              muxOutConnector[29] = fifoOut[34][9];
              muxOutConnector[30] = fifoOut[35][9];
              muxOutConnector[31] = fifoOut[36][9];
              muxOutConnector[32] = fifoOut[37][9];
              muxOutConnector[33] = fifoOut[38][9];
              muxOutConnector[34] = fifoOut[39][9];
              muxOutConnector[35] = fifoOut[40][9];
              muxOutConnector[36] = fifoOut[41][9];
              muxOutConnector[37] = fifoOut[42][9];
              muxOutConnector[38] = fifoOut[43][9];
              muxOutConnector[39] = fifoOut[44][9];
              muxOutConnector[40] = fifoOut[45][9];
              muxOutConnector[41] = fifoOut[46][9];
              muxOutConnector[42] = fifoOut[47][9];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
