`timescale 1ns / 1ps 
module InputQueueCirc_11(
        muxOut,
        rxIn,
        sliceAddress,
        wr_en,
        rd_en,
        clk,
        rst
);
parameter w = 6; // Width 
parameter maxVal = 63; // These are 0 LLRs 
parameter r = 32; // Rows of FIFO and input symbol count 
parameter c = 17; // Columns of FIFO
parameter muxOutSymbols = 52;
parameter ADDRESSWIDTH = 5;

parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 
output wire [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]rxIn;
input [ADDRESSWIDTH-1:0]sliceAddress;
input wr_en,rd_en;
 input clk,rst;

wire [ADDRESSWIDTH-1:0]sliceAddress_case;
wire [w-1:0]rxInConnector[r-1:0];
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output 
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign rxInConnector[k] = rxIn[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
           end  
        end
    end
    else if(wr_en) begin
        //LOAD inputs
            //Accept input
            for(i = r-1; i > -1; i=i-1) begin
               fifoOut[i][0] <= rxInConnector[i];
            end
        //Shifting process
        // Set (i,j)th value = (i,j-1)th value (except column 0)
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
    end
    else begin
       for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
       end
    end
end

assign sliceAddress_case = rd_en ? sliceAddress : READDISABLEDCASE;

// MUX WIRING
always@(*)begin
    case(sliceAddress_case)
       0: begin
              muxOutConnector[0] = fifoOut[21][16];
              muxOutConnector[1] = fifoOut[22][16];
              muxOutConnector[2] = fifoOut[23][16];
              muxOutConnector[3] = fifoOut[24][16];
              muxOutConnector[4] = fifoOut[25][16];
              muxOutConnector[5] = fifoOut[26][16];
              muxOutConnector[6] = fifoOut[27][16];
              muxOutConnector[7] = fifoOut[28][16];
              muxOutConnector[8] = fifoOut[29][16];
              muxOutConnector[9] = fifoOut[30][16];
              muxOutConnector[10] = fifoOut[31][16];
              muxOutConnector[11] = fifoOut[0][15];
              muxOutConnector[12] = fifoOut[1][15];
              muxOutConnector[13] = fifoOut[2][15];
              muxOutConnector[14] = fifoOut[3][15];
              muxOutConnector[15] = fifoOut[4][15];
              muxOutConnector[16] = fifoOut[5][15];
              muxOutConnector[17] = fifoOut[6][15];
              muxOutConnector[18] = fifoOut[7][15];
              muxOutConnector[19] = fifoOut[8][15];
              muxOutConnector[20] = fifoOut[9][15];
              muxOutConnector[21] = fifoOut[10][15];
              muxOutConnector[22] = fifoOut[11][15];
              muxOutConnector[23] = fifoOut[12][15];
              muxOutConnector[24] = fifoOut[13][15];
              muxOutConnector[25] = fifoOut[14][15];
              muxOutConnector[26] = fifoOut[28][8];
              muxOutConnector[27] = fifoOut[29][8];
              muxOutConnector[28] = fifoOut[30][8];
              muxOutConnector[29] = fifoOut[31][8];
              muxOutConnector[30] = fifoOut[0][7];
              muxOutConnector[31] = fifoOut[1][7];
              muxOutConnector[32] = fifoOut[2][7];
              muxOutConnector[33] = fifoOut[3][7];
              muxOutConnector[34] = fifoOut[4][7];
              muxOutConnector[35] = fifoOut[5][7];
              muxOutConnector[36] = fifoOut[6][7];
              muxOutConnector[37] = fifoOut[7][7];
              muxOutConnector[38] = fifoOut[8][7];
              muxOutConnector[39] = fifoOut[9][7];
              muxOutConnector[40] = fifoOut[10][7];
              muxOutConnector[41] = fifoOut[11][7];
              muxOutConnector[42] = fifoOut[12][7];
              muxOutConnector[43] = fifoOut[13][7];
              muxOutConnector[44] = fifoOut[14][7];
              muxOutConnector[45] = fifoOut[15][7];
              muxOutConnector[46] = fifoOut[16][7];
              muxOutConnector[47] = fifoOut[17][7];
              muxOutConnector[48] = fifoOut[18][7];
              muxOutConnector[49] = fifoOut[19][7];
              muxOutConnector[50] = fifoOut[20][7];
              muxOutConnector[51] = fifoOut[21][7];
       end
       1: begin
              muxOutConnector[0] = fifoOut[15][15];
              muxOutConnector[1] = fifoOut[16][15];
              muxOutConnector[2] = fifoOut[17][15];
              muxOutConnector[3] = fifoOut[18][15];
              muxOutConnector[4] = fifoOut[19][15];
              muxOutConnector[5] = fifoOut[20][15];
              muxOutConnector[6] = fifoOut[21][15];
              muxOutConnector[7] = fifoOut[22][15];
              muxOutConnector[8] = fifoOut[23][15];
              muxOutConnector[9] = fifoOut[24][15];
              muxOutConnector[10] = fifoOut[25][15];
              muxOutConnector[11] = fifoOut[26][15];
              muxOutConnector[12] = fifoOut[27][15];
              muxOutConnector[13] = fifoOut[28][15];
              muxOutConnector[14] = fifoOut[29][15];
              muxOutConnector[15] = fifoOut[30][15];
              muxOutConnector[16] = fifoOut[31][15];
              muxOutConnector[17] = fifoOut[0][14];
              muxOutConnector[18] = fifoOut[1][14];
              muxOutConnector[19] = fifoOut[2][14];
              muxOutConnector[20] = fifoOut[3][14];
              muxOutConnector[21] = fifoOut[4][14];
              muxOutConnector[22] = fifoOut[5][14];
              muxOutConnector[23] = fifoOut[6][14];
              muxOutConnector[24] = fifoOut[7][14];
              muxOutConnector[25] = fifoOut[8][14];
              muxOutConnector[26] = fifoOut[22][7];
              muxOutConnector[27] = fifoOut[23][7];
              muxOutConnector[28] = fifoOut[24][7];
              muxOutConnector[29] = fifoOut[25][7];
              muxOutConnector[30] = fifoOut[26][7];
              muxOutConnector[31] = fifoOut[27][7];
              muxOutConnector[32] = fifoOut[28][7];
              muxOutConnector[33] = fifoOut[29][7];
              muxOutConnector[34] = fifoOut[30][7];
              muxOutConnector[35] = fifoOut[31][7];
              muxOutConnector[36] = fifoOut[0][6];
              muxOutConnector[37] = fifoOut[1][6];
              muxOutConnector[38] = fifoOut[2][6];
              muxOutConnector[39] = fifoOut[3][6];
              muxOutConnector[40] = fifoOut[4][6];
              muxOutConnector[41] = fifoOut[5][6];
              muxOutConnector[42] = fifoOut[6][6];
              muxOutConnector[43] = fifoOut[7][6];
              muxOutConnector[44] = fifoOut[8][6];
              muxOutConnector[45] = fifoOut[9][6];
              muxOutConnector[46] = fifoOut[10][6];
              muxOutConnector[47] = fifoOut[11][6];
              muxOutConnector[48] = fifoOut[12][6];
              muxOutConnector[49] = fifoOut[13][6];
              muxOutConnector[50] = fifoOut[14][6];
              muxOutConnector[51] = fifoOut[15][6];
       end
       2: begin
              muxOutConnector[0] = fifoOut[9][14];
              muxOutConnector[1] = fifoOut[10][14];
              muxOutConnector[2] = fifoOut[11][14];
              muxOutConnector[3] = fifoOut[12][14];
              muxOutConnector[4] = fifoOut[13][14];
              muxOutConnector[5] = fifoOut[14][14];
              muxOutConnector[6] = fifoOut[15][14];
              muxOutConnector[7] = fifoOut[16][14];
              muxOutConnector[8] = fifoOut[17][14];
              muxOutConnector[9] = fifoOut[18][14];
              muxOutConnector[10] = fifoOut[19][14];
              muxOutConnector[11] = fifoOut[20][14];
              muxOutConnector[12] = fifoOut[21][14];
              muxOutConnector[13] = fifoOut[22][14];
              muxOutConnector[14] = fifoOut[23][14];
              muxOutConnector[15] = fifoOut[24][14];
              muxOutConnector[16] = fifoOut[25][14];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[0][13];
              muxOutConnector[24] = fifoOut[1][13];
              muxOutConnector[25] = fifoOut[2][13];
              muxOutConnector[26] = fifoOut[16][6];
              muxOutConnector[27] = fifoOut[17][6];
              muxOutConnector[28] = fifoOut[18][6];
              muxOutConnector[29] = fifoOut[19][6];
              muxOutConnector[30] = fifoOut[20][6];
              muxOutConnector[31] = fifoOut[21][6];
              muxOutConnector[32] = fifoOut[22][6];
              muxOutConnector[33] = fifoOut[23][6];
              muxOutConnector[34] = fifoOut[24][6];
              muxOutConnector[35] = fifoOut[25][6];
              muxOutConnector[36] = fifoOut[26][6];
              muxOutConnector[37] = fifoOut[27][6];
              muxOutConnector[38] = fifoOut[28][6];
              muxOutConnector[39] = fifoOut[29][6];
              muxOutConnector[40] = fifoOut[30][6];
              muxOutConnector[41] = fifoOut[31][6];
              muxOutConnector[42] = fifoOut[0][5];
              muxOutConnector[43] = fifoOut[1][5];
              muxOutConnector[44] = fifoOut[2][5];
              muxOutConnector[45] = fifoOut[3][5];
              muxOutConnector[46] = fifoOut[4][5];
              muxOutConnector[47] = fifoOut[5][5];
              muxOutConnector[48] = fifoOut[6][5];
              muxOutConnector[49] = fifoOut[7][5];
              muxOutConnector[50] = fifoOut[8][5];
              muxOutConnector[51] = fifoOut[9][5];
       end
       3: begin
              muxOutConnector[0] = fifoOut[3][13];
              muxOutConnector[1] = fifoOut[4][13];
              muxOutConnector[2] = fifoOut[5][13];
              muxOutConnector[3] = fifoOut[6][13];
              muxOutConnector[4] = fifoOut[7][13];
              muxOutConnector[5] = fifoOut[8][13];
              muxOutConnector[6] = fifoOut[9][13];
              muxOutConnector[7] = fifoOut[10][13];
              muxOutConnector[8] = fifoOut[11][13];
              muxOutConnector[9] = fifoOut[12][13];
              muxOutConnector[10] = fifoOut[13][13];
              muxOutConnector[11] = fifoOut[14][13];
              muxOutConnector[12] = fifoOut[15][13];
              muxOutConnector[13] = fifoOut[16][13];
              muxOutConnector[14] = fifoOut[17][13];
              muxOutConnector[15] = fifoOut[18][13];
              muxOutConnector[16] = fifoOut[19][13];
              muxOutConnector[17] = fifoOut[20][13];
              muxOutConnector[18] = fifoOut[21][13];
              muxOutConnector[19] = fifoOut[22][13];
              muxOutConnector[20] = fifoOut[23][13];
              muxOutConnector[21] = fifoOut[24][13];
              muxOutConnector[22] = fifoOut[25][13];
              muxOutConnector[23] = fifoOut[26][13];
              muxOutConnector[24] = fifoOut[27][13];
              muxOutConnector[25] = fifoOut[28][13];
              muxOutConnector[26] = fifoOut[10][5];
              muxOutConnector[27] = fifoOut[11][5];
              muxOutConnector[28] = fifoOut[12][5];
              muxOutConnector[29] = fifoOut[13][5];
              muxOutConnector[30] = fifoOut[14][5];
              muxOutConnector[31] = fifoOut[15][5];
              muxOutConnector[32] = fifoOut[16][5];
              muxOutConnector[33] = fifoOut[17][5];
              muxOutConnector[34] = fifoOut[18][5];
              muxOutConnector[35] = fifoOut[19][5];
              muxOutConnector[36] = fifoOut[20][5];
              muxOutConnector[37] = fifoOut[21][5];
              muxOutConnector[38] = fifoOut[22][5];
              muxOutConnector[39] = fifoOut[23][5];
              muxOutConnector[40] = fifoOut[24][5];
              muxOutConnector[41] = fifoOut[25][5];
              muxOutConnector[42] = fifoOut[26][5];
              muxOutConnector[43] = fifoOut[27][5];
              muxOutConnector[44] = fifoOut[28][5];
              muxOutConnector[45] = fifoOut[29][5];
              muxOutConnector[46] = fifoOut[30][5];
              muxOutConnector[47] = fifoOut[31][5];
              muxOutConnector[48] = fifoOut[0][4];
              muxOutConnector[49] = fifoOut[1][4];
              muxOutConnector[50] = fifoOut[2][4];
              muxOutConnector[51] = fifoOut[3][4];
       end
       4: begin
              muxOutConnector[0] = fifoOut[29][13];
              muxOutConnector[1] = fifoOut[30][13];
              muxOutConnector[2] = fifoOut[31][13];
              muxOutConnector[3] = fifoOut[0][12];
              muxOutConnector[4] = fifoOut[1][12];
              muxOutConnector[5] = fifoOut[2][12];
              muxOutConnector[6] = fifoOut[3][12];
              muxOutConnector[7] = fifoOut[4][12];
              muxOutConnector[8] = fifoOut[5][12];
              muxOutConnector[9] = fifoOut[6][12];
              muxOutConnector[10] = fifoOut[7][12];
              muxOutConnector[11] = fifoOut[8][12];
              muxOutConnector[12] = fifoOut[9][12];
              muxOutConnector[13] = fifoOut[10][12];
              muxOutConnector[14] = fifoOut[11][12];
              muxOutConnector[15] = fifoOut[12][12];
              muxOutConnector[16] = fifoOut[13][12];
              muxOutConnector[17] = fifoOut[14][12];
              muxOutConnector[18] = fifoOut[15][12];
              muxOutConnector[19] = fifoOut[16][12];
              muxOutConnector[20] = fifoOut[17][12];
              muxOutConnector[21] = fifoOut[18][12];
              muxOutConnector[22] = fifoOut[19][12];
              muxOutConnector[23] = fifoOut[20][12];
              muxOutConnector[24] = fifoOut[21][12];
              muxOutConnector[25] = fifoOut[22][12];
              muxOutConnector[26] = fifoOut[4][4];
              muxOutConnector[27] = fifoOut[5][4];
              muxOutConnector[28] = fifoOut[6][4];
              muxOutConnector[29] = fifoOut[7][4];
              muxOutConnector[30] = fifoOut[8][4];
              muxOutConnector[31] = fifoOut[9][4];
              muxOutConnector[32] = fifoOut[10][4];
              muxOutConnector[33] = fifoOut[11][4];
              muxOutConnector[34] = fifoOut[12][4];
              muxOutConnector[35] = fifoOut[13][4];
              muxOutConnector[36] = fifoOut[14][4];
              muxOutConnector[37] = fifoOut[15][4];
              muxOutConnector[38] = fifoOut[16][4];
              muxOutConnector[39] = fifoOut[17][4];
              muxOutConnector[40] = fifoOut[18][4];
              muxOutConnector[41] = fifoOut[19][4];
              muxOutConnector[42] = fifoOut[20][4];
              muxOutConnector[43] = fifoOut[21][4];
              muxOutConnector[44] = fifoOut[22][4];
              muxOutConnector[45] = fifoOut[23][4];
              muxOutConnector[46] = fifoOut[24][4];
              muxOutConnector[47] = fifoOut[25][4];
              muxOutConnector[48] = fifoOut[26][4];
              muxOutConnector[49] = fifoOut[27][4];
              muxOutConnector[50] = fifoOut[28][4];
              muxOutConnector[51] = fifoOut[29][4];
       end
       5: begin
              muxOutConnector[0] = fifoOut[23][12];
              muxOutConnector[1] = fifoOut[24][12];
              muxOutConnector[2] = fifoOut[25][12];
              muxOutConnector[3] = fifoOut[26][12];
              muxOutConnector[4] = fifoOut[27][12];
              muxOutConnector[5] = fifoOut[28][12];
              muxOutConnector[6] = fifoOut[29][12];
              muxOutConnector[7] = fifoOut[30][12];
              muxOutConnector[8] = fifoOut[31][12];
              muxOutConnector[9] = fifoOut[0][11];
              muxOutConnector[10] = fifoOut[1][11];
              muxOutConnector[11] = fifoOut[2][11];
              muxOutConnector[12] = fifoOut[3][11];
              muxOutConnector[13] = fifoOut[4][11];
              muxOutConnector[14] = fifoOut[5][11];
              muxOutConnector[15] = fifoOut[6][11];
              muxOutConnector[16] = fifoOut[7][11];
              muxOutConnector[17] = fifoOut[8][11];
              muxOutConnector[18] = fifoOut[9][11];
              muxOutConnector[19] = fifoOut[10][11];
              muxOutConnector[20] = fifoOut[11][11];
              muxOutConnector[21] = fifoOut[12][11];
              muxOutConnector[22] = fifoOut[13][11];
              muxOutConnector[23] = fifoOut[14][11];
              muxOutConnector[24] = fifoOut[15][11];
              muxOutConnector[25] = fifoOut[16][11];
              muxOutConnector[26] = fifoOut[30][4];
              muxOutConnector[27] = fifoOut[31][4];
              muxOutConnector[28] = fifoOut[0][3];
              muxOutConnector[29] = fifoOut[1][3];
              muxOutConnector[30] = fifoOut[2][3];
              muxOutConnector[31] = fifoOut[3][3];
              muxOutConnector[32] = fifoOut[4][3];
              muxOutConnector[33] = fifoOut[5][3];
              muxOutConnector[34] = fifoOut[6][3];
              muxOutConnector[35] = fifoOut[7][3];
              muxOutConnector[36] = fifoOut[8][3];
              muxOutConnector[37] = fifoOut[9][3];
              muxOutConnector[38] = fifoOut[10][3];
              muxOutConnector[39] = fifoOut[11][3];
              muxOutConnector[40] = fifoOut[12][3];
              muxOutConnector[41] = fifoOut[13][3];
              muxOutConnector[42] = fifoOut[14][3];
              muxOutConnector[43] = fifoOut[15][3];
              muxOutConnector[44] = fifoOut[16][3];
              muxOutConnector[45] = fifoOut[17][3];
              muxOutConnector[46] = fifoOut[18][3];
              muxOutConnector[47] = fifoOut[19][3];
              muxOutConnector[48] = fifoOut[20][3];
              muxOutConnector[49] = fifoOut[21][3];
              muxOutConnector[50] = fifoOut[22][3];
              muxOutConnector[51] = fifoOut[23][3];
       end
       6: begin
              muxOutConnector[0] = fifoOut[17][11];
              muxOutConnector[1] = fifoOut[18][11];
              muxOutConnector[2] = fifoOut[19][11];
              muxOutConnector[3] = fifoOut[20][11];
              muxOutConnector[4] = fifoOut[21][11];
              muxOutConnector[5] = fifoOut[22][11];
              muxOutConnector[6] = fifoOut[23][11];
              muxOutConnector[7] = fifoOut[24][11];
              muxOutConnector[8] = fifoOut[25][11];
              muxOutConnector[9] = fifoOut[26][11];
              muxOutConnector[10] = fifoOut[27][11];
              muxOutConnector[11] = fifoOut[28][11];
              muxOutConnector[12] = fifoOut[29][11];
              muxOutConnector[13] = fifoOut[30][11];
              muxOutConnector[14] = fifoOut[31][11];
              muxOutConnector[15] = fifoOut[0][10];
              muxOutConnector[16] = fifoOut[1][10];
              muxOutConnector[17] = fifoOut[2][10];
              muxOutConnector[18] = fifoOut[3][10];
              muxOutConnector[19] = fifoOut[4][10];
              muxOutConnector[20] = fifoOut[5][10];
              muxOutConnector[21] = fifoOut[6][10];
              muxOutConnector[22] = fifoOut[7][10];
              muxOutConnector[23] = fifoOut[8][10];
              muxOutConnector[24] = fifoOut[9][10];
              muxOutConnector[25] = fifoOut[10][10];
              muxOutConnector[26] = fifoOut[24][3];
              muxOutConnector[27] = fifoOut[25][3];
              muxOutConnector[28] = fifoOut[26][3];
              muxOutConnector[29] = fifoOut[27][3];
              muxOutConnector[30] = fifoOut[28][3];
              muxOutConnector[31] = fifoOut[29][3];
              muxOutConnector[32] = fifoOut[30][3];
              muxOutConnector[33] = fifoOut[31][3];
              muxOutConnector[34] = fifoOut[0][2];
              muxOutConnector[35] = fifoOut[1][2];
              muxOutConnector[36] = fifoOut[2][2];
              muxOutConnector[37] = fifoOut[3][2];
              muxOutConnector[38] = fifoOut[4][2];
              muxOutConnector[39] = fifoOut[5][2];
              muxOutConnector[40] = fifoOut[6][2];
              muxOutConnector[41] = fifoOut[7][2];
              muxOutConnector[42] = fifoOut[8][2];
              muxOutConnector[43] = fifoOut[9][2];
              muxOutConnector[44] = fifoOut[10][2];
              muxOutConnector[45] = fifoOut[11][2];
              muxOutConnector[46] = fifoOut[12][2];
              muxOutConnector[47] = fifoOut[13][2];
              muxOutConnector[48] = fifoOut[14][2];
              muxOutConnector[49] = fifoOut[15][2];
              muxOutConnector[50] = fifoOut[16][2];
              muxOutConnector[51] = fifoOut[17][2];
       end
       7: begin
              muxOutConnector[0] = fifoOut[11][10];
              muxOutConnector[1] = fifoOut[12][10];
              muxOutConnector[2] = fifoOut[13][10];
              muxOutConnector[3] = fifoOut[14][10];
              muxOutConnector[4] = fifoOut[15][10];
              muxOutConnector[5] = fifoOut[16][10];
              muxOutConnector[6] = fifoOut[17][10];
              muxOutConnector[7] = fifoOut[18][10];
              muxOutConnector[8] = fifoOut[19][10];
              muxOutConnector[9] = fifoOut[20][10];
              muxOutConnector[10] = fifoOut[21][10];
              muxOutConnector[11] = fifoOut[22][10];
              muxOutConnector[12] = fifoOut[23][10];
              muxOutConnector[13] = fifoOut[24][10];
              muxOutConnector[14] = fifoOut[25][10];
              muxOutConnector[15] = fifoOut[26][10];
              muxOutConnector[16] = fifoOut[27][10];
              muxOutConnector[17] = fifoOut[28][10];
              muxOutConnector[18] = fifoOut[29][10];
              muxOutConnector[19] = fifoOut[30][10];
              muxOutConnector[20] = fifoOut[31][10];
              muxOutConnector[21] = fifoOut[0][9];
              muxOutConnector[22] = fifoOut[1][9];
              muxOutConnector[23] = fifoOut[2][9];
              muxOutConnector[24] = fifoOut[3][9];
              muxOutConnector[25] = fifoOut[4][9];
              muxOutConnector[26] = fifoOut[18][2];
              muxOutConnector[27] = fifoOut[19][2];
              muxOutConnector[28] = fifoOut[20][2];
              muxOutConnector[29] = fifoOut[21][2];
              muxOutConnector[30] = fifoOut[22][2];
              muxOutConnector[31] = fifoOut[23][2];
              muxOutConnector[32] = fifoOut[24][2];
              muxOutConnector[33] = fifoOut[25][2];
              muxOutConnector[34] = fifoOut[26][2];
              muxOutConnector[35] = fifoOut[27][2];
              muxOutConnector[36] = fifoOut[28][2];
              muxOutConnector[37] = fifoOut[29][2];
              muxOutConnector[38] = fifoOut[30][2];
              muxOutConnector[39] = fifoOut[31][2];
              muxOutConnector[40] = fifoOut[0][1];
              muxOutConnector[41] = fifoOut[1][1];
              muxOutConnector[42] = fifoOut[2][1];
              muxOutConnector[43] = fifoOut[3][1];
              muxOutConnector[44] = fifoOut[4][1];
              muxOutConnector[45] = fifoOut[5][1];
              muxOutConnector[46] = fifoOut[6][1];
              muxOutConnector[47] = fifoOut[7][1];
              muxOutConnector[48] = fifoOut[8][1];
              muxOutConnector[49] = fifoOut[9][1];
              muxOutConnector[50] = fifoOut[10][1];
              muxOutConnector[51] = fifoOut[11][1];
       end
       8: begin
              muxOutConnector[0] = fifoOut[5][9];
              muxOutConnector[1] = fifoOut[6][9];
              muxOutConnector[2] = fifoOut[7][9];
              muxOutConnector[3] = fifoOut[8][9];
              muxOutConnector[4] = fifoOut[9][9];
              muxOutConnector[5] = fifoOut[10][9];
              muxOutConnector[6] = fifoOut[11][9];
              muxOutConnector[7] = fifoOut[12][9];
              muxOutConnector[8] = fifoOut[13][9];
              muxOutConnector[9] = fifoOut[14][9];
              muxOutConnector[10] = fifoOut[15][9];
              muxOutConnector[11] = fifoOut[16][9];
              muxOutConnector[12] = fifoOut[17][9];
              muxOutConnector[13] = fifoOut[18][9];
              muxOutConnector[14] = fifoOut[19][9];
              muxOutConnector[15] = fifoOut[20][9];
              muxOutConnector[16] = fifoOut[21][9];
              muxOutConnector[17] = fifoOut[22][9];
              muxOutConnector[18] = fifoOut[23][9];
              muxOutConnector[19] = fifoOut[24][9];
              muxOutConnector[20] = fifoOut[25][9];
              muxOutConnector[21] = fifoOut[26][9];
              muxOutConnector[22] = fifoOut[27][9];
              muxOutConnector[23] = fifoOut[28][9];
              muxOutConnector[24] = fifoOut[29][9];
              muxOutConnector[25] = fifoOut[30][9];
              muxOutConnector[26] = fifoOut[12][1];
              muxOutConnector[27] = fifoOut[13][1];
              muxOutConnector[28] = fifoOut[14][1];
              muxOutConnector[29] = fifoOut[15][1];
              muxOutConnector[30] = fifoOut[16][1];
              muxOutConnector[31] = fifoOut[17][1];
              muxOutConnector[32] = fifoOut[18][1];
              muxOutConnector[33] = fifoOut[19][1];
              muxOutConnector[34] = fifoOut[20][1];
              muxOutConnector[35] = fifoOut[21][1];
              muxOutConnector[36] = fifoOut[22][1];
              muxOutConnector[37] = fifoOut[23][1];
              muxOutConnector[38] = fifoOut[24][1];
              muxOutConnector[39] = fifoOut[25][1];
              muxOutConnector[40] = fifoOut[26][1];
              muxOutConnector[41] = fifoOut[27][1];
              muxOutConnector[42] = fifoOut[28][1];
              muxOutConnector[43] = fifoOut[29][1];
              muxOutConnector[44] = fifoOut[30][1];
              muxOutConnector[45] = fifoOut[31][1];
              muxOutConnector[46] = fifoOut[0][0];
              muxOutConnector[47] = fifoOut[1][0];
              muxOutConnector[48] = fifoOut[3][16];
              muxOutConnector[49] = fifoOut[4][16];
              muxOutConnector[50] = fifoOut[5][16];
              muxOutConnector[51] = fifoOut[6][16];
       end
       9: begin
              muxOutConnector[0] = fifoOut[31][9];
              muxOutConnector[1] = fifoOut[0][8];
              muxOutConnector[2] = fifoOut[1][8];
              muxOutConnector[3] = fifoOut[2][8];
              muxOutConnector[4] = fifoOut[3][8];
              muxOutConnector[5] = fifoOut[4][8];
              muxOutConnector[6] = fifoOut[5][8];
              muxOutConnector[7] = fifoOut[6][8];
              muxOutConnector[8] = fifoOut[7][8];
              muxOutConnector[9] = fifoOut[8][8];
              muxOutConnector[10] = fifoOut[9][8];
              muxOutConnector[11] = fifoOut[10][8];
              muxOutConnector[12] = fifoOut[11][8];
              muxOutConnector[13] = fifoOut[12][8];
              muxOutConnector[14] = fifoOut[13][8];
              muxOutConnector[15] = fifoOut[14][8];
              muxOutConnector[16] = fifoOut[15][8];
              muxOutConnector[17] = fifoOut[16][8];
              muxOutConnector[18] = fifoOut[17][8];
              muxOutConnector[19] = fifoOut[18][8];
              muxOutConnector[20] = fifoOut[19][8];
              muxOutConnector[21] = fifoOut[20][8];
              muxOutConnector[22] = fifoOut[21][8];
              muxOutConnector[23] = fifoOut[22][8];
              muxOutConnector[24] = fifoOut[23][8];
              muxOutConnector[25] = fifoOut[24][8];
              muxOutConnector[26] = fifoOut[7][16];
              muxOutConnector[27] = fifoOut[8][16];
              muxOutConnector[28] = fifoOut[9][16];
              muxOutConnector[29] = fifoOut[10][16];
              muxOutConnector[30] = fifoOut[11][16];
              muxOutConnector[31] = fifoOut[12][16];
              muxOutConnector[32] = fifoOut[13][16];
              muxOutConnector[33] = fifoOut[14][16];
              muxOutConnector[34] = fifoOut[15][16];
              muxOutConnector[35] = fifoOut[16][16];
              muxOutConnector[36] = fifoOut[17][16];
              muxOutConnector[37] = fifoOut[18][16];
              muxOutConnector[38] = fifoOut[19][16];
              muxOutConnector[39] = fifoOut[20][16];
              muxOutConnector[40] = fifoOut[21][16];
              muxOutConnector[41] = fifoOut[22][16];
              muxOutConnector[42] = fifoOut[23][16];
              muxOutConnector[43] = fifoOut[24][16];
              muxOutConnector[44] = fifoOut[25][16];
              muxOutConnector[45] = fifoOut[26][16];
              muxOutConnector[46] = fifoOut[27][16];
              muxOutConnector[47] = fifoOut[28][16];
              muxOutConnector[48] = fifoOut[29][16];
              muxOutConnector[49] = fifoOut[30][16];
              muxOutConnector[50] = fifoOut[31][16];
              muxOutConnector[51] = fifoOut[0][15];
       end
       10: begin
              muxOutConnector[0] = fifoOut[25][8];
              muxOutConnector[1] = fifoOut[26][8];
              muxOutConnector[2] = fifoOut[27][8];
              muxOutConnector[3] = fifoOut[28][8];
              muxOutConnector[4] = fifoOut[29][8];
              muxOutConnector[5] = fifoOut[30][8];
              muxOutConnector[6] = fifoOut[31][8];
              muxOutConnector[7] = fifoOut[0][7];
              muxOutConnector[8] = fifoOut[1][7];
              muxOutConnector[9] = fifoOut[2][7];
              muxOutConnector[10] = fifoOut[3][7];
              muxOutConnector[11] = fifoOut[4][7];
              muxOutConnector[12] = fifoOut[5][7];
              muxOutConnector[13] = fifoOut[6][7];
              muxOutConnector[14] = fifoOut[7][7];
              muxOutConnector[15] = fifoOut[8][7];
              muxOutConnector[16] = fifoOut[9][7];
              muxOutConnector[17] = fifoOut[10][7];
              muxOutConnector[18] = fifoOut[11][7];
              muxOutConnector[19] = fifoOut[12][7];
              muxOutConnector[20] = fifoOut[13][7];
              muxOutConnector[21] = fifoOut[14][7];
              muxOutConnector[22] = fifoOut[15][7];
              muxOutConnector[23] = fifoOut[16][7];
              muxOutConnector[24] = fifoOut[17][7];
              muxOutConnector[25] = fifoOut[18][7];
              muxOutConnector[26] = fifoOut[1][15];
              muxOutConnector[27] = fifoOut[2][15];
              muxOutConnector[28] = fifoOut[3][15];
              muxOutConnector[29] = fifoOut[4][15];
              muxOutConnector[30] = fifoOut[5][15];
              muxOutConnector[31] = fifoOut[6][15];
              muxOutConnector[32] = fifoOut[7][15];
              muxOutConnector[33] = fifoOut[8][15];
              muxOutConnector[34] = fifoOut[9][15];
              muxOutConnector[35] = fifoOut[10][15];
              muxOutConnector[36] = fifoOut[11][15];
              muxOutConnector[37] = fifoOut[12][15];
              muxOutConnector[38] = fifoOut[13][15];
              muxOutConnector[39] = fifoOut[14][15];
              muxOutConnector[40] = fifoOut[15][15];
              muxOutConnector[41] = fifoOut[16][15];
              muxOutConnector[42] = fifoOut[17][15];
              muxOutConnector[43] = fifoOut[18][15];
              muxOutConnector[44] = fifoOut[19][15];
              muxOutConnector[45] = fifoOut[20][15];
              muxOutConnector[46] = fifoOut[21][15];
              muxOutConnector[47] = fifoOut[22][15];
              muxOutConnector[48] = fifoOut[23][15];
              muxOutConnector[49] = fifoOut[24][15];
              muxOutConnector[50] = fifoOut[25][15];
              muxOutConnector[51] = fifoOut[26][15];
       end
       11: begin
              muxOutConnector[0] = fifoOut[19][7];
              muxOutConnector[1] = fifoOut[20][7];
              muxOutConnector[2] = fifoOut[21][7];
              muxOutConnector[3] = fifoOut[22][7];
              muxOutConnector[4] = fifoOut[23][7];
              muxOutConnector[5] = fifoOut[24][7];
              muxOutConnector[6] = fifoOut[25][7];
              muxOutConnector[7] = fifoOut[26][7];
              muxOutConnector[8] = fifoOut[27][7];
              muxOutConnector[9] = fifoOut[28][7];
              muxOutConnector[10] = fifoOut[29][7];
              muxOutConnector[11] = fifoOut[30][7];
              muxOutConnector[12] = fifoOut[31][7];
              muxOutConnector[13] = fifoOut[0][6];
              muxOutConnector[14] = fifoOut[1][6];
              muxOutConnector[15] = fifoOut[2][6];
              muxOutConnector[16] = fifoOut[3][6];
              muxOutConnector[17] = fifoOut[4][6];
              muxOutConnector[18] = fifoOut[5][6];
              muxOutConnector[19] = fifoOut[6][6];
              muxOutConnector[20] = fifoOut[7][6];
              muxOutConnector[21] = fifoOut[8][6];
              muxOutConnector[22] = fifoOut[9][6];
              muxOutConnector[23] = fifoOut[10][6];
              muxOutConnector[24] = fifoOut[11][6];
              muxOutConnector[25] = fifoOut[12][6];
              muxOutConnector[26] = fifoOut[27][15];
              muxOutConnector[27] = fifoOut[28][15];
              muxOutConnector[28] = fifoOut[29][15];
              muxOutConnector[29] = fifoOut[30][15];
              muxOutConnector[30] = fifoOut[31][15];
              muxOutConnector[31] = fifoOut[0][14];
              muxOutConnector[32] = fifoOut[1][14];
              muxOutConnector[33] = fifoOut[2][14];
              muxOutConnector[34] = fifoOut[3][14];
              muxOutConnector[35] = fifoOut[4][14];
              muxOutConnector[36] = fifoOut[5][14];
              muxOutConnector[37] = fifoOut[6][14];
              muxOutConnector[38] = fifoOut[7][14];
              muxOutConnector[39] = fifoOut[8][14];
              muxOutConnector[40] = fifoOut[9][14];
              muxOutConnector[41] = fifoOut[10][14];
              muxOutConnector[42] = fifoOut[11][14];
              muxOutConnector[43] = fifoOut[12][14];
              muxOutConnector[44] = fifoOut[13][14];
              muxOutConnector[45] = fifoOut[14][14];
              muxOutConnector[46] = fifoOut[15][14];
              muxOutConnector[47] = fifoOut[16][14];
              muxOutConnector[48] = fifoOut[17][14];
              muxOutConnector[49] = fifoOut[18][14];
              muxOutConnector[50] = fifoOut[19][14];
              muxOutConnector[51] = fifoOut[20][14];
       end
       12: begin
              muxOutConnector[0] = fifoOut[13][6];
              muxOutConnector[1] = fifoOut[14][6];
              muxOutConnector[2] = fifoOut[15][6];
              muxOutConnector[3] = fifoOut[16][6];
              muxOutConnector[4] = fifoOut[17][6];
              muxOutConnector[5] = fifoOut[18][6];
              muxOutConnector[6] = fifoOut[19][6];
              muxOutConnector[7] = fifoOut[20][6];
              muxOutConnector[8] = fifoOut[21][6];
              muxOutConnector[9] = fifoOut[22][6];
              muxOutConnector[10] = fifoOut[23][6];
              muxOutConnector[11] = fifoOut[24][6];
              muxOutConnector[12] = fifoOut[25][6];
              muxOutConnector[13] = fifoOut[26][6];
              muxOutConnector[14] = fifoOut[27][6];
              muxOutConnector[15] = fifoOut[28][6];
              muxOutConnector[16] = fifoOut[29][6];
              muxOutConnector[17] = fifoOut[30][6];
              muxOutConnector[18] = fifoOut[31][6];
              muxOutConnector[19] = fifoOut[0][5];
              muxOutConnector[20] = fifoOut[1][5];
              muxOutConnector[21] = fifoOut[2][5];
              muxOutConnector[22] = fifoOut[3][5];
              muxOutConnector[23] = fifoOut[4][5];
              muxOutConnector[24] = fifoOut[5][5];
              muxOutConnector[25] = fifoOut[6][5];
              muxOutConnector[26] = fifoOut[21][14];
              muxOutConnector[27] = fifoOut[22][14];
              muxOutConnector[28] = fifoOut[23][14];
              muxOutConnector[29] = fifoOut[24][14];
              muxOutConnector[30] = fifoOut[25][14];
              muxOutConnector[31] = fifoOut[26][14];
              muxOutConnector[32] = fifoOut[27][14];
              muxOutConnector[33] = fifoOut[28][14];
              muxOutConnector[34] = fifoOut[29][14];
              muxOutConnector[35] = fifoOut[30][14];
              muxOutConnector[36] = fifoOut[31][14];
              muxOutConnector[37] = fifoOut[0][13];
              muxOutConnector[38] = fifoOut[1][13];
              muxOutConnector[39] = fifoOut[2][13];
              muxOutConnector[40] = fifoOut[3][13];
              muxOutConnector[41] = fifoOut[4][13];
              muxOutConnector[42] = fifoOut[5][13];
              muxOutConnector[43] = fifoOut[6][13];
              muxOutConnector[44] = fifoOut[7][13];
              muxOutConnector[45] = fifoOut[8][13];
              muxOutConnector[46] = fifoOut[9][13];
              muxOutConnector[47] = fifoOut[10][13];
              muxOutConnector[48] = fifoOut[11][13];
              muxOutConnector[49] = fifoOut[12][13];
              muxOutConnector[50] = fifoOut[13][13];
              muxOutConnector[51] = fifoOut[14][13];
       end
       13: begin
              muxOutConnector[0] = fifoOut[7][5];
              muxOutConnector[1] = fifoOut[8][5];
              muxOutConnector[2] = fifoOut[9][5];
              muxOutConnector[3] = fifoOut[10][5];
              muxOutConnector[4] = fifoOut[11][5];
              muxOutConnector[5] = fifoOut[12][5];
              muxOutConnector[6] = fifoOut[13][5];
              muxOutConnector[7] = fifoOut[14][5];
              muxOutConnector[8] = fifoOut[15][5];
              muxOutConnector[9] = fifoOut[16][5];
              muxOutConnector[10] = fifoOut[17][5];
              muxOutConnector[11] = fifoOut[18][5];
              muxOutConnector[12] = fifoOut[19][5];
              muxOutConnector[13] = fifoOut[20][5];
              muxOutConnector[14] = fifoOut[21][5];
              muxOutConnector[15] = fifoOut[22][5];
              muxOutConnector[16] = fifoOut[23][5];
              muxOutConnector[17] = fifoOut[24][5];
              muxOutConnector[18] = fifoOut[25][5];
              muxOutConnector[19] = fifoOut[26][5];
              muxOutConnector[20] = fifoOut[27][5];
              muxOutConnector[21] = fifoOut[28][5];
              muxOutConnector[22] = fifoOut[29][5];
              muxOutConnector[23] = fifoOut[30][5];
              muxOutConnector[24] = fifoOut[31][5];
              muxOutConnector[25] = fifoOut[0][4];
              muxOutConnector[26] = fifoOut[15][13];
              muxOutConnector[27] = fifoOut[16][13];
              muxOutConnector[28] = fifoOut[17][13];
              muxOutConnector[29] = fifoOut[18][13];
              muxOutConnector[30] = fifoOut[19][13];
              muxOutConnector[31] = fifoOut[20][13];
              muxOutConnector[32] = fifoOut[21][13];
              muxOutConnector[33] = fifoOut[22][13];
              muxOutConnector[34] = fifoOut[23][13];
              muxOutConnector[35] = fifoOut[24][13];
              muxOutConnector[36] = fifoOut[25][13];
              muxOutConnector[37] = fifoOut[26][13];
              muxOutConnector[38] = fifoOut[27][13];
              muxOutConnector[39] = fifoOut[28][13];
              muxOutConnector[40] = fifoOut[29][13];
              muxOutConnector[41] = fifoOut[30][13];
              muxOutConnector[42] = fifoOut[31][13];
              muxOutConnector[43] = fifoOut[0][12];
              muxOutConnector[44] = fifoOut[1][12];
              muxOutConnector[45] = fifoOut[2][12];
              muxOutConnector[46] = fifoOut[3][12];
              muxOutConnector[47] = fifoOut[4][12];
              muxOutConnector[48] = fifoOut[5][12];
              muxOutConnector[49] = fifoOut[6][12];
              muxOutConnector[50] = fifoOut[7][12];
              muxOutConnector[51] = fifoOut[8][12];
       end
       14: begin
              muxOutConnector[0] = fifoOut[1][4];
              muxOutConnector[1] = fifoOut[2][4];
              muxOutConnector[2] = fifoOut[3][4];
              muxOutConnector[3] = fifoOut[4][4];
              muxOutConnector[4] = fifoOut[5][4];
              muxOutConnector[5] = fifoOut[6][4];
              muxOutConnector[6] = fifoOut[7][4];
              muxOutConnector[7] = fifoOut[8][4];
              muxOutConnector[8] = fifoOut[9][4];
              muxOutConnector[9] = fifoOut[10][4];
              muxOutConnector[10] = fifoOut[11][4];
              muxOutConnector[11] = fifoOut[12][4];
              muxOutConnector[12] = fifoOut[13][4];
              muxOutConnector[13] = fifoOut[14][4];
              muxOutConnector[14] = fifoOut[15][4];
              muxOutConnector[15] = fifoOut[16][4];
              muxOutConnector[16] = fifoOut[17][4];
              muxOutConnector[17] = fifoOut[18][4];
              muxOutConnector[18] = fifoOut[19][4];
              muxOutConnector[19] = fifoOut[20][4];
              muxOutConnector[20] = fifoOut[21][4];
              muxOutConnector[21] = fifoOut[22][4];
              muxOutConnector[22] = fifoOut[23][4];
              muxOutConnector[23] = fifoOut[24][4];
              muxOutConnector[24] = fifoOut[25][4];
              muxOutConnector[25] = fifoOut[26][4];
              muxOutConnector[26] = fifoOut[9][12];
              muxOutConnector[27] = fifoOut[10][12];
              muxOutConnector[28] = fifoOut[11][12];
              muxOutConnector[29] = fifoOut[12][12];
              muxOutConnector[30] = fifoOut[13][12];
              muxOutConnector[31] = fifoOut[14][12];
              muxOutConnector[32] = fifoOut[15][12];
              muxOutConnector[33] = fifoOut[16][12];
              muxOutConnector[34] = fifoOut[17][12];
              muxOutConnector[35] = fifoOut[18][12];
              muxOutConnector[36] = fifoOut[19][12];
              muxOutConnector[37] = fifoOut[20][12];
              muxOutConnector[38] = fifoOut[21][12];
              muxOutConnector[39] = fifoOut[22][12];
              muxOutConnector[40] = fifoOut[23][12];
              muxOutConnector[41] = fifoOut[24][12];
              muxOutConnector[42] = fifoOut[25][12];
              muxOutConnector[43] = fifoOut[26][12];
              muxOutConnector[44] = fifoOut[27][12];
              muxOutConnector[45] = fifoOut[28][12];
              muxOutConnector[46] = fifoOut[29][12];
              muxOutConnector[47] = fifoOut[30][12];
              muxOutConnector[48] = fifoOut[31][12];
              muxOutConnector[49] = fifoOut[0][11];
              muxOutConnector[50] = fifoOut[1][11];
              muxOutConnector[51] = fifoOut[2][11];
       end
       15: begin
              muxOutConnector[0] = fifoOut[27][4];
              muxOutConnector[1] = fifoOut[28][4];
              muxOutConnector[2] = fifoOut[29][4];
              muxOutConnector[3] = fifoOut[30][4];
              muxOutConnector[4] = fifoOut[31][4];
              muxOutConnector[5] = fifoOut[0][3];
              muxOutConnector[6] = fifoOut[1][3];
              muxOutConnector[7] = fifoOut[2][3];
              muxOutConnector[8] = fifoOut[3][3];
              muxOutConnector[9] = fifoOut[4][3];
              muxOutConnector[10] = fifoOut[5][3];
              muxOutConnector[11] = fifoOut[6][3];
              muxOutConnector[12] = fifoOut[7][3];
              muxOutConnector[13] = fifoOut[8][3];
              muxOutConnector[14] = fifoOut[9][3];
              muxOutConnector[15] = fifoOut[10][3];
              muxOutConnector[16] = fifoOut[11][3];
              muxOutConnector[17] = fifoOut[12][3];
              muxOutConnector[18] = fifoOut[13][3];
              muxOutConnector[19] = fifoOut[14][3];
              muxOutConnector[20] = fifoOut[15][3];
              muxOutConnector[21] = fifoOut[16][3];
              muxOutConnector[22] = fifoOut[17][3];
              muxOutConnector[23] = fifoOut[18][3];
              muxOutConnector[24] = fifoOut[19][3];
              muxOutConnector[25] = fifoOut[20][3];
              muxOutConnector[26] = fifoOut[3][11];
              muxOutConnector[27] = fifoOut[4][11];
              muxOutConnector[28] = fifoOut[5][11];
              muxOutConnector[29] = fifoOut[6][11];
              muxOutConnector[30] = fifoOut[7][11];
              muxOutConnector[31] = fifoOut[8][11];
              muxOutConnector[32] = fifoOut[9][11];
              muxOutConnector[33] = fifoOut[10][11];
              muxOutConnector[34] = fifoOut[11][11];
              muxOutConnector[35] = fifoOut[12][11];
              muxOutConnector[36] = fifoOut[13][11];
              muxOutConnector[37] = fifoOut[14][11];
              muxOutConnector[38] = fifoOut[15][11];
              muxOutConnector[39] = fifoOut[16][11];
              muxOutConnector[40] = fifoOut[17][11];
              muxOutConnector[41] = fifoOut[18][11];
              muxOutConnector[42] = fifoOut[19][11];
              muxOutConnector[43] = fifoOut[20][11];
              muxOutConnector[44] = fifoOut[21][11];
              muxOutConnector[45] = fifoOut[22][11];
              muxOutConnector[46] = fifoOut[23][11];
              muxOutConnector[47] = fifoOut[24][11];
              muxOutConnector[48] = fifoOut[25][11];
              muxOutConnector[49] = fifoOut[26][11];
              muxOutConnector[50] = fifoOut[27][11];
              muxOutConnector[51] = fifoOut[28][11];
       end
       16: begin
              muxOutConnector[0] = fifoOut[21][3];
              muxOutConnector[1] = fifoOut[22][3];
              muxOutConnector[2] = fifoOut[23][3];
              muxOutConnector[3] = fifoOut[24][3];
              muxOutConnector[4] = fifoOut[25][3];
              muxOutConnector[5] = fifoOut[26][3];
              muxOutConnector[6] = fifoOut[27][3];
              muxOutConnector[7] = fifoOut[28][3];
              muxOutConnector[8] = fifoOut[29][3];
              muxOutConnector[9] = fifoOut[30][3];
              muxOutConnector[10] = fifoOut[31][3];
              muxOutConnector[11] = fifoOut[0][2];
              muxOutConnector[12] = fifoOut[1][2];
              muxOutConnector[13] = fifoOut[2][2];
              muxOutConnector[14] = fifoOut[3][2];
              muxOutConnector[15] = fifoOut[4][2];
              muxOutConnector[16] = fifoOut[5][2];
              muxOutConnector[17] = fifoOut[6][2];
              muxOutConnector[18] = fifoOut[7][2];
              muxOutConnector[19] = fifoOut[8][2];
              muxOutConnector[20] = fifoOut[9][2];
              muxOutConnector[21] = fifoOut[10][2];
              muxOutConnector[22] = fifoOut[11][2];
              muxOutConnector[23] = fifoOut[12][2];
              muxOutConnector[24] = fifoOut[13][2];
              muxOutConnector[25] = fifoOut[14][2];
              muxOutConnector[26] = fifoOut[29][11];
              muxOutConnector[27] = fifoOut[30][11];
              muxOutConnector[28] = fifoOut[31][11];
              muxOutConnector[29] = fifoOut[0][10];
              muxOutConnector[30] = fifoOut[1][10];
              muxOutConnector[31] = fifoOut[2][10];
              muxOutConnector[32] = fifoOut[3][10];
              muxOutConnector[33] = fifoOut[4][10];
              muxOutConnector[34] = fifoOut[5][10];
              muxOutConnector[35] = fifoOut[6][10];
              muxOutConnector[36] = fifoOut[7][10];
              muxOutConnector[37] = fifoOut[8][10];
              muxOutConnector[38] = fifoOut[9][10];
              muxOutConnector[39] = fifoOut[10][10];
              muxOutConnector[40] = fifoOut[11][10];
              muxOutConnector[41] = fifoOut[12][10];
              muxOutConnector[42] = fifoOut[13][10];
              muxOutConnector[43] = fifoOut[14][10];
              muxOutConnector[44] = fifoOut[15][10];
              muxOutConnector[45] = fifoOut[16][10];
              muxOutConnector[46] = fifoOut[17][10];
              muxOutConnector[47] = fifoOut[18][10];
              muxOutConnector[48] = fifoOut[19][10];
              muxOutConnector[49] = fifoOut[20][10];
              muxOutConnector[50] = fifoOut[21][10];
              muxOutConnector[51] = fifoOut[22][10];
       end
       17: begin
              muxOutConnector[0] = fifoOut[15][2];
              muxOutConnector[1] = fifoOut[16][2];
              muxOutConnector[2] = fifoOut[17][2];
              muxOutConnector[3] = fifoOut[18][2];
              muxOutConnector[4] = fifoOut[19][2];
              muxOutConnector[5] = fifoOut[20][2];
              muxOutConnector[6] = fifoOut[21][2];
              muxOutConnector[7] = fifoOut[22][2];
              muxOutConnector[8] = fifoOut[23][2];
              muxOutConnector[9] = fifoOut[24][2];
              muxOutConnector[10] = fifoOut[25][2];
              muxOutConnector[11] = fifoOut[26][2];
              muxOutConnector[12] = fifoOut[27][2];
              muxOutConnector[13] = fifoOut[28][2];
              muxOutConnector[14] = fifoOut[29][2];
              muxOutConnector[15] = fifoOut[30][2];
              muxOutConnector[16] = fifoOut[31][2];
              muxOutConnector[17] = fifoOut[0][1];
              muxOutConnector[18] = fifoOut[1][1];
              muxOutConnector[19] = fifoOut[2][1];
              muxOutConnector[20] = fifoOut[3][1];
              muxOutConnector[21] = fifoOut[4][1];
              muxOutConnector[22] = fifoOut[5][1];
              muxOutConnector[23] = fifoOut[6][1];
              muxOutConnector[24] = fifoOut[7][1];
              muxOutConnector[25] = fifoOut[8][1];
              muxOutConnector[26] = fifoOut[23][10];
              muxOutConnector[27] = fifoOut[24][10];
              muxOutConnector[28] = fifoOut[25][10];
              muxOutConnector[29] = fifoOut[26][10];
              muxOutConnector[30] = fifoOut[27][10];
              muxOutConnector[31] = fifoOut[28][10];
              muxOutConnector[32] = fifoOut[29][10];
              muxOutConnector[33] = fifoOut[30][10];
              muxOutConnector[34] = fifoOut[31][10];
              muxOutConnector[35] = fifoOut[0][9];
              muxOutConnector[36] = fifoOut[1][9];
              muxOutConnector[37] = fifoOut[2][9];
              muxOutConnector[38] = fifoOut[3][9];
              muxOutConnector[39] = fifoOut[4][9];
              muxOutConnector[40] = fifoOut[5][9];
              muxOutConnector[41] = fifoOut[6][9];
              muxOutConnector[42] = fifoOut[7][9];
              muxOutConnector[43] = fifoOut[8][9];
              muxOutConnector[44] = fifoOut[9][9];
              muxOutConnector[45] = fifoOut[10][9];
              muxOutConnector[46] = fifoOut[11][9];
              muxOutConnector[47] = fifoOut[12][9];
              muxOutConnector[48] = fifoOut[13][9];
              muxOutConnector[49] = fifoOut[14][9];
              muxOutConnector[50] = fifoOut[15][9];
              muxOutConnector[51] = fifoOut[16][9];
       end
       18: begin
              muxOutConnector[0] = fifoOut[9][1];
              muxOutConnector[1] = fifoOut[10][1];
              muxOutConnector[2] = fifoOut[11][1];
              muxOutConnector[3] = fifoOut[12][1];
              muxOutConnector[4] = fifoOut[13][1];
              muxOutConnector[5] = fifoOut[14][1];
              muxOutConnector[6] = fifoOut[15][1];
              muxOutConnector[7] = fifoOut[16][1];
              muxOutConnector[8] = fifoOut[17][1];
              muxOutConnector[9] = fifoOut[18][1];
              muxOutConnector[10] = fifoOut[19][1];
              muxOutConnector[11] = fifoOut[20][1];
              muxOutConnector[12] = fifoOut[21][1];
              muxOutConnector[13] = fifoOut[22][1];
              muxOutConnector[14] = fifoOut[23][1];
              muxOutConnector[15] = fifoOut[24][1];
              muxOutConnector[16] = fifoOut[25][1];
              muxOutConnector[17] = fifoOut[26][1];
              muxOutConnector[18] = fifoOut[27][1];
              muxOutConnector[19] = fifoOut[28][1];
              muxOutConnector[20] = fifoOut[29][1];
              muxOutConnector[21] = fifoOut[30][1];
              muxOutConnector[22] = fifoOut[31][1];
              muxOutConnector[23] = fifoOut[0][0];
              muxOutConnector[24] = fifoOut[1][0];
              muxOutConnector[25] = fifoOut[3][16];
              muxOutConnector[26] = fifoOut[17][9];
              muxOutConnector[27] = fifoOut[18][9];
              muxOutConnector[28] = fifoOut[19][9];
              muxOutConnector[29] = fifoOut[20][9];
              muxOutConnector[30] = fifoOut[21][9];
              muxOutConnector[31] = fifoOut[22][9];
              muxOutConnector[32] = fifoOut[23][9];
              muxOutConnector[33] = fifoOut[24][9];
              muxOutConnector[34] = fifoOut[25][9];
              muxOutConnector[35] = fifoOut[26][9];
              muxOutConnector[36] = fifoOut[27][9];
              muxOutConnector[37] = fifoOut[28][9];
              muxOutConnector[38] = fifoOut[29][9];
              muxOutConnector[39] = fifoOut[30][9];
              muxOutConnector[40] = fifoOut[31][9];
              muxOutConnector[41] = fifoOut[0][8];
              muxOutConnector[42] = fifoOut[1][8];
              muxOutConnector[43] = fifoOut[2][8];
              muxOutConnector[44] = fifoOut[3][8];
              muxOutConnector[45] = fifoOut[4][8];
              muxOutConnector[46] = fifoOut[5][8];
              muxOutConnector[47] = fifoOut[6][8];
              muxOutConnector[48] = fifoOut[7][8];
              muxOutConnector[49] = fifoOut[8][8];
              muxOutConnector[50] = fifoOut[9][8];
              muxOutConnector[51] = fifoOut[10][8];
       end
       19: begin
              muxOutConnector[0] = fifoOut[4][16];
              muxOutConnector[1] = fifoOut[5][16];
              muxOutConnector[2] = fifoOut[6][16];
              muxOutConnector[3] = fifoOut[7][16];
              muxOutConnector[4] = fifoOut[8][16];
              muxOutConnector[5] = fifoOut[9][16];
              muxOutConnector[6] = fifoOut[10][16];
              muxOutConnector[7] = fifoOut[11][16];
              muxOutConnector[8] = fifoOut[12][16];
              muxOutConnector[9] = fifoOut[13][16];
              muxOutConnector[10] = fifoOut[14][16];
              muxOutConnector[11] = fifoOut[15][16];
              muxOutConnector[12] = fifoOut[16][16];
              muxOutConnector[13] = fifoOut[17][16];
              muxOutConnector[14] = fifoOut[18][16];
              muxOutConnector[15] = fifoOut[19][16];
              muxOutConnector[16] = fifoOut[20][16];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[11][8];
              muxOutConnector[27] = fifoOut[12][8];
              muxOutConnector[28] = fifoOut[13][8];
              muxOutConnector[29] = fifoOut[14][8];
              muxOutConnector[30] = fifoOut[15][8];
              muxOutConnector[31] = fifoOut[16][8];
              muxOutConnector[32] = fifoOut[17][8];
              muxOutConnector[33] = fifoOut[18][8];
              muxOutConnector[34] = fifoOut[19][8];
              muxOutConnector[35] = fifoOut[20][8];
              muxOutConnector[36] = fifoOut[21][8];
              muxOutConnector[37] = fifoOut[22][8];
              muxOutConnector[38] = fifoOut[23][8];
              muxOutConnector[39] = fifoOut[24][8];
              muxOutConnector[40] = fifoOut[25][8];
              muxOutConnector[41] = fifoOut[26][8];
              muxOutConnector[42] = fifoOut[27][8];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
