`timescale 1ns / 1ps
module LMem1To0_511_circ10_combined_ys_yu_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        rxIn,
        load_input_en,
        iteration_0_indicator,
        feedback_en,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter r_lower = 32;
parameter c = 17;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input load_input_en;
input iteration_0_indicator;
input [ADDRESSWIDTH-1:0]unloadAddress;
input feedback_en;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input [ r_lower * w - 1 : 0 ] rxIn; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
wire [w-1:0]rxInConnector[r_lower-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

generate
    for (k=0;k<r_lower;k=k+1)begin:assign_rx
        assign rxInConnector[k] = rxIn[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            if(feedback_en)begin
                 fifoOut[i][0] <= fifoOut[i][c-1];
            end
            else if(load_input_en)begin
                 if(i < r_lower)begin
                   fifoOut[i][0] = rxInConnector[i];
                 end
                 else begin
                   fifoOut[i][0] = maxVal;
                 end
            end
            else begin
                 fifoOut[i][0] <= ly0InConnector[i];
            end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
       0: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = fifoOut[25][4][w-1];
              unloadMuxOut[23] = fifoOut[0][3][w-1];
              unloadMuxOut[24] = fifoOut[1][3][w-1];
              unloadMuxOut[25] = fifoOut[2][3][w-1];
              unloadMuxOut[26] = fifoOut[3][3][w-1];
              unloadMuxOut[27] = fifoOut[4][3][w-1];
              unloadMuxOut[28] = fifoOut[5][3][w-1];
              unloadMuxOut[29] = fifoOut[6][3][w-1];
              unloadMuxOut[30] = fifoOut[7][3][w-1];
              unloadMuxOut[31] = fifoOut[8][3][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[9][4][w-1];
              unloadMuxOut[1] = fifoOut[10][4][w-1];
              unloadMuxOut[2] = fifoOut[11][4][w-1];
              unloadMuxOut[3] = fifoOut[12][4][w-1];
              unloadMuxOut[4] = fifoOut[13][4][w-1];
              unloadMuxOut[5] = fifoOut[14][4][w-1];
              unloadMuxOut[6] = fifoOut[15][4][w-1];
              unloadMuxOut[7] = fifoOut[16][4][w-1];
              unloadMuxOut[8] = fifoOut[17][4][w-1];
              unloadMuxOut[9] = fifoOut[18][4][w-1];
              unloadMuxOut[10] = fifoOut[19][4][w-1];
              unloadMuxOut[11] = fifoOut[20][4][w-1];
              unloadMuxOut[12] = fifoOut[21][4][w-1];
              unloadMuxOut[13] = fifoOut[22][4][w-1];
              unloadMuxOut[14] = fifoOut[23][4][w-1];
              unloadMuxOut[15] = fifoOut[24][4][w-1];
              unloadMuxOut[16] = fifoOut[25][4][w-1];
              unloadMuxOut[17] = fifoOut[0][3][w-1];
              unloadMuxOut[18] = fifoOut[1][3][w-1];
              unloadMuxOut[19] = fifoOut[2][3][w-1];
              unloadMuxOut[20] = fifoOut[3][3][w-1];
              unloadMuxOut[21] = fifoOut[4][3][w-1];
              unloadMuxOut[22] = fifoOut[5][3][w-1];
              unloadMuxOut[23] = fifoOut[6][3][w-1];
              unloadMuxOut[24] = fifoOut[7][3][w-1];
              unloadMuxOut[25] = fifoOut[8][3][w-1];
              unloadMuxOut[26] = fifoOut[9][3][w-1];
              unloadMuxOut[27] = fifoOut[10][3][w-1];
              unloadMuxOut[28] = fifoOut[11][3][w-1];
              unloadMuxOut[29] = fifoOut[12][3][w-1];
              unloadMuxOut[30] = fifoOut[13][3][w-1];
              unloadMuxOut[31] = fifoOut[14][3][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[15][4][w-1];
              unloadMuxOut[1] = fifoOut[16][4][w-1];
              unloadMuxOut[2] = fifoOut[17][4][w-1];
              unloadMuxOut[3] = fifoOut[18][4][w-1];
              unloadMuxOut[4] = fifoOut[19][4][w-1];
              unloadMuxOut[5] = fifoOut[20][4][w-1];
              unloadMuxOut[6] = fifoOut[21][4][w-1];
              unloadMuxOut[7] = fifoOut[22][4][w-1];
              unloadMuxOut[8] = fifoOut[23][4][w-1];
              unloadMuxOut[9] = fifoOut[24][4][w-1];
              unloadMuxOut[10] = fifoOut[25][4][w-1];
              unloadMuxOut[11] = fifoOut[0][3][w-1];
              unloadMuxOut[12] = fifoOut[1][3][w-1];
              unloadMuxOut[13] = fifoOut[2][3][w-1];
              unloadMuxOut[14] = fifoOut[3][3][w-1];
              unloadMuxOut[15] = fifoOut[4][3][w-1];
              unloadMuxOut[16] = fifoOut[5][3][w-1];
              unloadMuxOut[17] = fifoOut[6][3][w-1];
              unloadMuxOut[18] = fifoOut[7][3][w-1];
              unloadMuxOut[19] = fifoOut[8][3][w-1];
              unloadMuxOut[20] = fifoOut[9][3][w-1];
              unloadMuxOut[21] = fifoOut[10][3][w-1];
              unloadMuxOut[22] = fifoOut[11][3][w-1];
              unloadMuxOut[23] = fifoOut[12][3][w-1];
              unloadMuxOut[24] = fifoOut[13][3][w-1];
              unloadMuxOut[25] = fifoOut[14][3][w-1];
              unloadMuxOut[26] = fifoOut[15][3][w-1];
              unloadMuxOut[27] = fifoOut[16][3][w-1];
              unloadMuxOut[28] = fifoOut[17][3][w-1];
              unloadMuxOut[29] = fifoOut[18][3][w-1];
              unloadMuxOut[30] = fifoOut[19][3][w-1];
              unloadMuxOut[31] = fifoOut[20][3][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[21][4][w-1];
              unloadMuxOut[1] = fifoOut[22][4][w-1];
              unloadMuxOut[2] = fifoOut[26][14][w-1];
              unloadMuxOut[3] = fifoOut[27][14][w-1];
              unloadMuxOut[4] = fifoOut[28][14][w-1];
              unloadMuxOut[5] = fifoOut[29][14][w-1];
              unloadMuxOut[6] = fifoOut[30][14][w-1];
              unloadMuxOut[7] = fifoOut[31][14][w-1];
              unloadMuxOut[8] = fifoOut[32][14][w-1];
              unloadMuxOut[9] = fifoOut[33][14][w-1];
              unloadMuxOut[10] = fifoOut[34][14][w-1];
              unloadMuxOut[11] = fifoOut[35][14][w-1];
              unloadMuxOut[12] = fifoOut[36][14][w-1];
              unloadMuxOut[13] = fifoOut[37][14][w-1];
              unloadMuxOut[14] = fifoOut[38][14][w-1];
              unloadMuxOut[15] = fifoOut[39][14][w-1];
              unloadMuxOut[16] = fifoOut[40][14][w-1];
              unloadMuxOut[17] = fifoOut[41][14][w-1];
              unloadMuxOut[18] = fifoOut[42][14][w-1];
              unloadMuxOut[19] = fifoOut[43][14][w-1];
              unloadMuxOut[20] = fifoOut[44][14][w-1];
              unloadMuxOut[21] = fifoOut[45][14][w-1];
              unloadMuxOut[22] = fifoOut[46][14][w-1];
              unloadMuxOut[23] = fifoOut[47][14][w-1];
              unloadMuxOut[24] = fifoOut[48][14][w-1];
              unloadMuxOut[25] = fifoOut[49][14][w-1];
              unloadMuxOut[26] = fifoOut[50][14][w-1];
              unloadMuxOut[27] = fifoOut[51][14][w-1];
              unloadMuxOut[28] = fifoOut[26][13][w-1];
              unloadMuxOut[29] = fifoOut[27][13][w-1];
              unloadMuxOut[30] = fifoOut[28][13][w-1];
              unloadMuxOut[31] = fifoOut[29][13][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[30][14][w-1];
              unloadMuxOut[1] = fifoOut[31][14][w-1];
              unloadMuxOut[2] = fifoOut[32][14][w-1];
              unloadMuxOut[3] = fifoOut[33][14][w-1];
              unloadMuxOut[4] = fifoOut[34][14][w-1];
              unloadMuxOut[5] = fifoOut[35][14][w-1];
              unloadMuxOut[6] = fifoOut[36][14][w-1];
              unloadMuxOut[7] = fifoOut[37][14][w-1];
              unloadMuxOut[8] = fifoOut[38][14][w-1];
              unloadMuxOut[9] = fifoOut[39][14][w-1];
              unloadMuxOut[10] = fifoOut[40][14][w-1];
              unloadMuxOut[11] = fifoOut[41][14][w-1];
              unloadMuxOut[12] = fifoOut[42][14][w-1];
              unloadMuxOut[13] = fifoOut[43][14][w-1];
              unloadMuxOut[14] = fifoOut[44][14][w-1];
              unloadMuxOut[15] = fifoOut[45][14][w-1];
              unloadMuxOut[16] = fifoOut[46][14][w-1];
              unloadMuxOut[17] = fifoOut[47][14][w-1];
              unloadMuxOut[18] = fifoOut[48][14][w-1];
              unloadMuxOut[19] = fifoOut[49][14][w-1];
              unloadMuxOut[20] = fifoOut[50][14][w-1];
              unloadMuxOut[21] = fifoOut[51][14][w-1];
              unloadMuxOut[22] = fifoOut[26][13][w-1];
              unloadMuxOut[23] = fifoOut[27][13][w-1];
              unloadMuxOut[24] = fifoOut[28][13][w-1];
              unloadMuxOut[25] = fifoOut[29][13][w-1];
              unloadMuxOut[26] = fifoOut[30][13][w-1];
              unloadMuxOut[27] = fifoOut[31][13][w-1];
              unloadMuxOut[28] = fifoOut[32][13][w-1];
              unloadMuxOut[29] = fifoOut[33][13][w-1];
              unloadMuxOut[30] = fifoOut[34][13][w-1];
              unloadMuxOut[31] = fifoOut[35][13][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[36][14][w-1];
              unloadMuxOut[1] = fifoOut[37][14][w-1];
              unloadMuxOut[2] = fifoOut[38][14][w-1];
              unloadMuxOut[3] = fifoOut[39][14][w-1];
              unloadMuxOut[4] = fifoOut[40][14][w-1];
              unloadMuxOut[5] = fifoOut[41][14][w-1];
              unloadMuxOut[6] = fifoOut[42][14][w-1];
              unloadMuxOut[7] = fifoOut[43][14][w-1];
              unloadMuxOut[8] = fifoOut[44][14][w-1];
              unloadMuxOut[9] = fifoOut[45][14][w-1];
              unloadMuxOut[10] = fifoOut[46][14][w-1];
              unloadMuxOut[11] = fifoOut[47][14][w-1];
              unloadMuxOut[12] = fifoOut[48][14][w-1];
              unloadMuxOut[13] = fifoOut[49][14][w-1];
              unloadMuxOut[14] = fifoOut[50][14][w-1];
              unloadMuxOut[15] = fifoOut[51][14][w-1];
              unloadMuxOut[16] = fifoOut[26][13][w-1];
              unloadMuxOut[17] = fifoOut[27][13][w-1];
              unloadMuxOut[18] = fifoOut[28][13][w-1];
              unloadMuxOut[19] = fifoOut[29][13][w-1];
              unloadMuxOut[20] = fifoOut[30][13][w-1];
              unloadMuxOut[21] = fifoOut[31][13][w-1];
              unloadMuxOut[22] = fifoOut[32][13][w-1];
              unloadMuxOut[23] = fifoOut[33][13][w-1];
              unloadMuxOut[24] = fifoOut[34][13][w-1];
              unloadMuxOut[25] = fifoOut[35][13][w-1];
              unloadMuxOut[26] = fifoOut[36][13][w-1];
              unloadMuxOut[27] = fifoOut[37][13][w-1];
              unloadMuxOut[28] = fifoOut[38][13][w-1];
              unloadMuxOut[29] = fifoOut[39][13][w-1];
              unloadMuxOut[30] = fifoOut[40][13][w-1];
              unloadMuxOut[31] = fifoOut[41][13][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[42][14][w-1];
              unloadMuxOut[1] = fifoOut[43][14][w-1];
              unloadMuxOut[2] = fifoOut[44][14][w-1];
              unloadMuxOut[3] = fifoOut[45][14][w-1];
              unloadMuxOut[4] = fifoOut[46][14][w-1];
              unloadMuxOut[5] = fifoOut[47][14][w-1];
              unloadMuxOut[6] = fifoOut[48][14][w-1];
              unloadMuxOut[7] = fifoOut[49][14][w-1];
              unloadMuxOut[8] = fifoOut[50][14][w-1];
              unloadMuxOut[9] = fifoOut[51][14][w-1];
              unloadMuxOut[10] = fifoOut[26][13][w-1];
              unloadMuxOut[11] = fifoOut[27][13][w-1];
              unloadMuxOut[12] = fifoOut[28][13][w-1];
              unloadMuxOut[13] = fifoOut[29][13][w-1];
              unloadMuxOut[14] = fifoOut[30][13][w-1];
              unloadMuxOut[15] = fifoOut[31][13][w-1];
              unloadMuxOut[16] = fifoOut[32][13][w-1];
              unloadMuxOut[17] = fifoOut[33][13][w-1];
              unloadMuxOut[18] = fifoOut[34][13][w-1];
              unloadMuxOut[19] = fifoOut[35][13][w-1];
              unloadMuxOut[20] = fifoOut[36][13][w-1];
              unloadMuxOut[21] = fifoOut[37][13][w-1];
              unloadMuxOut[22] = fifoOut[38][13][w-1];
              unloadMuxOut[23] = fifoOut[39][13][w-1];
              unloadMuxOut[24] = fifoOut[40][13][w-1];
              unloadMuxOut[25] = fifoOut[41][13][w-1];
              unloadMuxOut[26] = fifoOut[42][13][w-1];
              unloadMuxOut[27] = fifoOut[43][13][w-1];
              unloadMuxOut[28] = fifoOut[44][13][w-1];
              unloadMuxOut[29] = fifoOut[45][13][w-1];
              unloadMuxOut[30] = fifoOut[46][13][w-1];
              unloadMuxOut[31] = fifoOut[47][13][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[48][14][w-1];
              unloadMuxOut[1] = fifoOut[49][14][w-1];
              unloadMuxOut[2] = fifoOut[50][14][w-1];
              unloadMuxOut[3] = fifoOut[51][14][w-1];
              unloadMuxOut[4] = fifoOut[26][13][w-1];
              unloadMuxOut[5] = fifoOut[27][13][w-1];
              unloadMuxOut[6] = fifoOut[28][13][w-1];
              unloadMuxOut[7] = fifoOut[29][13][w-1];
              unloadMuxOut[8] = fifoOut[30][13][w-1];
              unloadMuxOut[9] = fifoOut[31][13][w-1];
              unloadMuxOut[10] = fifoOut[32][13][w-1];
              unloadMuxOut[11] = fifoOut[33][13][w-1];
              unloadMuxOut[12] = fifoOut[34][13][w-1];
              unloadMuxOut[13] = fifoOut[35][13][w-1];
              unloadMuxOut[14] = fifoOut[36][13][w-1];
              unloadMuxOut[15] = fifoOut[37][13][w-1];
              unloadMuxOut[16] = fifoOut[38][13][w-1];
              unloadMuxOut[17] = fifoOut[39][13][w-1];
              unloadMuxOut[18] = fifoOut[40][13][w-1];
              unloadMuxOut[19] = fifoOut[41][13][w-1];
              unloadMuxOut[20] = fifoOut[42][13][w-1];
              unloadMuxOut[21] = fifoOut[43][13][w-1];
              unloadMuxOut[22] = fifoOut[44][13][w-1];
              unloadMuxOut[23] = fifoOut[45][13][w-1];
              unloadMuxOut[24] = fifoOut[46][13][w-1];
              unloadMuxOut[25] = fifoOut[47][13][w-1];
              unloadMuxOut[26] = fifoOut[48][13][w-1];
              unloadMuxOut[27] = fifoOut[49][13][w-1];
              unloadMuxOut[28] = fifoOut[50][13][w-1];
              unloadMuxOut[29] = fifoOut[51][13][w-1];
              unloadMuxOut[30] = fifoOut[26][12][w-1];
              unloadMuxOut[31] = fifoOut[27][12][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[28][13][w-1];
              unloadMuxOut[1] = fifoOut[29][13][w-1];
              unloadMuxOut[2] = fifoOut[30][13][w-1];
              unloadMuxOut[3] = fifoOut[31][13][w-1];
              unloadMuxOut[4] = fifoOut[32][13][w-1];
              unloadMuxOut[5] = fifoOut[33][13][w-1];
              unloadMuxOut[6] = fifoOut[34][13][w-1];
              unloadMuxOut[7] = fifoOut[35][13][w-1];
              unloadMuxOut[8] = fifoOut[36][13][w-1];
              unloadMuxOut[9] = fifoOut[37][13][w-1];
              unloadMuxOut[10] = fifoOut[38][13][w-1];
              unloadMuxOut[11] = fifoOut[39][13][w-1];
              unloadMuxOut[12] = fifoOut[40][13][w-1];
              unloadMuxOut[13] = fifoOut[41][13][w-1];
              unloadMuxOut[14] = fifoOut[42][13][w-1];
              unloadMuxOut[15] = fifoOut[43][13][w-1];
              unloadMuxOut[16] = fifoOut[44][13][w-1];
              unloadMuxOut[17] = fifoOut[45][13][w-1];
              unloadMuxOut[18] = fifoOut[46][13][w-1];
              unloadMuxOut[19] = fifoOut[47][13][w-1];
              unloadMuxOut[20] = fifoOut[48][13][w-1];
              unloadMuxOut[21] = fifoOut[49][13][w-1];
              unloadMuxOut[22] = fifoOut[50][13][w-1];
              unloadMuxOut[23] = fifoOut[51][13][w-1];
              unloadMuxOut[24] = fifoOut[26][12][w-1];
              unloadMuxOut[25] = fifoOut[27][12][w-1];
              unloadMuxOut[26] = fifoOut[28][12][w-1];
              unloadMuxOut[27] = fifoOut[29][12][w-1];
              unloadMuxOut[28] = fifoOut[30][12][w-1];
              unloadMuxOut[29] = fifoOut[31][12][w-1];
              unloadMuxOut[30] = fifoOut[32][12][w-1];
              unloadMuxOut[31] = fifoOut[33][12][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[34][13][w-1];
              unloadMuxOut[1] = fifoOut[35][13][w-1];
              unloadMuxOut[2] = fifoOut[36][13][w-1];
              unloadMuxOut[3] = fifoOut[37][13][w-1];
              unloadMuxOut[4] = fifoOut[38][13][w-1];
              unloadMuxOut[5] = fifoOut[39][13][w-1];
              unloadMuxOut[6] = fifoOut[40][13][w-1];
              unloadMuxOut[7] = fifoOut[41][13][w-1];
              unloadMuxOut[8] = fifoOut[42][13][w-1];
              unloadMuxOut[9] = fifoOut[43][13][w-1];
              unloadMuxOut[10] = fifoOut[44][13][w-1];
              unloadMuxOut[11] = fifoOut[45][13][w-1];
              unloadMuxOut[12] = fifoOut[46][13][w-1];
              unloadMuxOut[13] = fifoOut[47][13][w-1];
              unloadMuxOut[14] = fifoOut[48][13][w-1];
              unloadMuxOut[15] = fifoOut[49][13][w-1];
              unloadMuxOut[16] = fifoOut[50][13][w-1];
              unloadMuxOut[17] = fifoOut[51][13][w-1];
              unloadMuxOut[18] = fifoOut[26][12][w-1];
              unloadMuxOut[19] = fifoOut[27][12][w-1];
              unloadMuxOut[20] = fifoOut[28][12][w-1];
              unloadMuxOut[21] = fifoOut[29][12][w-1];
              unloadMuxOut[22] = fifoOut[30][12][w-1];
              unloadMuxOut[23] = fifoOut[31][12][w-1];
              unloadMuxOut[24] = fifoOut[32][12][w-1];
              unloadMuxOut[25] = fifoOut[33][12][w-1];
              unloadMuxOut[26] = fifoOut[34][12][w-1];
              unloadMuxOut[27] = fifoOut[35][12][w-1];
              unloadMuxOut[28] = fifoOut[36][12][w-1];
              unloadMuxOut[29] = fifoOut[37][12][w-1];
              unloadMuxOut[30] = fifoOut[38][12][w-1];
              unloadMuxOut[31] = fifoOut[39][12][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[40][13][w-1];
              unloadMuxOut[1] = fifoOut[41][13][w-1];
              unloadMuxOut[2] = fifoOut[42][13][w-1];
              unloadMuxOut[3] = fifoOut[43][13][w-1];
              unloadMuxOut[4] = fifoOut[44][13][w-1];
              unloadMuxOut[5] = fifoOut[45][13][w-1];
              unloadMuxOut[6] = fifoOut[46][13][w-1];
              unloadMuxOut[7] = fifoOut[47][13][w-1];
              unloadMuxOut[8] = fifoOut[48][13][w-1];
              unloadMuxOut[9] = fifoOut[49][13][w-1];
              unloadMuxOut[10] = fifoOut[50][13][w-1];
              unloadMuxOut[11] = fifoOut[51][13][w-1];
              unloadMuxOut[12] = fifoOut[26][12][w-1];
              unloadMuxOut[13] = fifoOut[27][12][w-1];
              unloadMuxOut[14] = fifoOut[28][12][w-1];
              unloadMuxOut[15] = fifoOut[29][12][w-1];
              unloadMuxOut[16] = fifoOut[30][12][w-1];
              unloadMuxOut[17] = fifoOut[31][12][w-1];
              unloadMuxOut[18] = fifoOut[32][12][w-1];
              unloadMuxOut[19] = fifoOut[33][12][w-1];
              unloadMuxOut[20] = fifoOut[34][12][w-1];
              unloadMuxOut[21] = fifoOut[35][12][w-1];
              unloadMuxOut[22] = fifoOut[36][12][w-1];
              unloadMuxOut[23] = fifoOut[37][12][w-1];
              unloadMuxOut[24] = fifoOut[38][12][w-1];
              unloadMuxOut[25] = fifoOut[39][12][w-1];
              unloadMuxOut[26] = fifoOut[40][12][w-1];
              unloadMuxOut[27] = fifoOut[41][12][w-1];
              unloadMuxOut[28] = fifoOut[42][12][w-1];
              unloadMuxOut[29] = fifoOut[43][12][w-1];
              unloadMuxOut[30] = fifoOut[44][12][w-1];
              unloadMuxOut[31] = fifoOut[45][12][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[46][13][w-1];
              unloadMuxOut[1] = fifoOut[47][13][w-1];
              unloadMuxOut[2] = fifoOut[48][13][w-1];
              unloadMuxOut[3] = fifoOut[49][13][w-1];
              unloadMuxOut[4] = fifoOut[50][13][w-1];
              unloadMuxOut[5] = fifoOut[51][13][w-1];
              unloadMuxOut[6] = fifoOut[26][12][w-1];
              unloadMuxOut[7] = fifoOut[27][12][w-1];
              unloadMuxOut[8] = fifoOut[28][12][w-1];
              unloadMuxOut[9] = fifoOut[29][12][w-1];
              unloadMuxOut[10] = fifoOut[30][12][w-1];
              unloadMuxOut[11] = fifoOut[31][12][w-1];
              unloadMuxOut[12] = fifoOut[32][12][w-1];
              unloadMuxOut[13] = fifoOut[33][12][w-1];
              unloadMuxOut[14] = fifoOut[34][12][w-1];
              unloadMuxOut[15] = fifoOut[35][12][w-1];
              unloadMuxOut[16] = fifoOut[36][12][w-1];
              unloadMuxOut[17] = fifoOut[37][12][w-1];
              unloadMuxOut[18] = fifoOut[38][12][w-1];
              unloadMuxOut[19] = fifoOut[39][12][w-1];
              unloadMuxOut[20] = fifoOut[40][12][w-1];
              unloadMuxOut[21] = fifoOut[41][12][w-1];
              unloadMuxOut[22] = fifoOut[42][12][w-1];
              unloadMuxOut[23] = fifoOut[43][12][w-1];
              unloadMuxOut[24] = fifoOut[44][12][w-1];
              unloadMuxOut[25] = fifoOut[45][12][w-1];
              unloadMuxOut[26] = fifoOut[46][12][w-1];
              unloadMuxOut[27] = fifoOut[47][12][w-1];
              unloadMuxOut[28] = fifoOut[48][12][w-1];
              unloadMuxOut[29] = fifoOut[49][12][w-1];
              unloadMuxOut[30] = fifoOut[50][12][w-1];
              unloadMuxOut[31] = fifoOut[51][12][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[26][12][w-1];
              unloadMuxOut[1] = fifoOut[27][12][w-1];
              unloadMuxOut[2] = fifoOut[28][12][w-1];
              unloadMuxOut[3] = fifoOut[29][12][w-1];
              unloadMuxOut[4] = fifoOut[30][12][w-1];
              unloadMuxOut[5] = fifoOut[31][12][w-1];
              unloadMuxOut[6] = fifoOut[32][12][w-1];
              unloadMuxOut[7] = fifoOut[33][12][w-1];
              unloadMuxOut[8] = fifoOut[34][12][w-1];
              unloadMuxOut[9] = fifoOut[35][12][w-1];
              unloadMuxOut[10] = fifoOut[36][12][w-1];
              unloadMuxOut[11] = fifoOut[37][12][w-1];
              unloadMuxOut[12] = fifoOut[38][12][w-1];
              unloadMuxOut[13] = fifoOut[39][12][w-1];
              unloadMuxOut[14] = fifoOut[40][12][w-1];
              unloadMuxOut[15] = fifoOut[41][12][w-1];
              unloadMuxOut[16] = fifoOut[42][12][w-1];
              unloadMuxOut[17] = fifoOut[23][4][w-1];
              unloadMuxOut[18] = fifoOut[24][4][w-1];
              unloadMuxOut[19] = fifoOut[25][4][w-1];
              unloadMuxOut[20] = fifoOut[0][3][w-1];
              unloadMuxOut[21] = fifoOut[1][3][w-1];
              unloadMuxOut[22] = fifoOut[2][3][w-1];
              unloadMuxOut[23] = fifoOut[3][3][w-1];
              unloadMuxOut[24] = fifoOut[4][3][w-1];
              unloadMuxOut[25] = fifoOut[5][3][w-1];
              unloadMuxOut[26] = fifoOut[6][3][w-1];
              unloadMuxOut[27] = fifoOut[7][3][w-1];
              unloadMuxOut[28] = fifoOut[8][3][w-1];
              unloadMuxOut[29] = fifoOut[9][3][w-1];
              unloadMuxOut[30] = fifoOut[10][3][w-1];
              unloadMuxOut[31] = fifoOut[11][3][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[12][4][w-1];
              unloadMuxOut[1] = fifoOut[13][4][w-1];
              unloadMuxOut[2] = fifoOut[14][4][w-1];
              unloadMuxOut[3] = fifoOut[15][4][w-1];
              unloadMuxOut[4] = fifoOut[16][4][w-1];
              unloadMuxOut[5] = fifoOut[17][4][w-1];
              unloadMuxOut[6] = fifoOut[18][4][w-1];
              unloadMuxOut[7] = fifoOut[19][4][w-1];
              unloadMuxOut[8] = fifoOut[20][4][w-1];
              unloadMuxOut[9] = fifoOut[21][4][w-1];
              unloadMuxOut[10] = fifoOut[22][4][w-1];
              unloadMuxOut[11] = fifoOut[23][4][w-1];
              unloadMuxOut[12] = fifoOut[24][4][w-1];
              unloadMuxOut[13] = fifoOut[25][4][w-1];
              unloadMuxOut[14] = fifoOut[0][3][w-1];
              unloadMuxOut[15] = fifoOut[1][3][w-1];
              unloadMuxOut[16] = fifoOut[2][3][w-1];
              unloadMuxOut[17] = fifoOut[3][3][w-1];
              unloadMuxOut[18] = fifoOut[4][3][w-1];
              unloadMuxOut[19] = fifoOut[5][3][w-1];
              unloadMuxOut[20] = fifoOut[6][3][w-1];
              unloadMuxOut[21] = fifoOut[7][3][w-1];
              unloadMuxOut[22] = fifoOut[8][3][w-1];
              unloadMuxOut[23] = fifoOut[9][3][w-1];
              unloadMuxOut[24] = fifoOut[10][3][w-1];
              unloadMuxOut[25] = fifoOut[11][3][w-1];
              unloadMuxOut[26] = fifoOut[12][3][w-1];
              unloadMuxOut[27] = fifoOut[13][3][w-1];
              unloadMuxOut[28] = fifoOut[14][3][w-1];
              unloadMuxOut[29] = fifoOut[15][3][w-1];
              unloadMuxOut[30] = fifoOut[16][3][w-1];
              unloadMuxOut[31] = fifoOut[17][3][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[18][4][w-1];
              unloadMuxOut[1] = fifoOut[19][4][w-1];
              unloadMuxOut[2] = fifoOut[20][4][w-1];
              unloadMuxOut[3] = fifoOut[21][4][w-1];
              unloadMuxOut[4] = fifoOut[22][4][w-1];
              unloadMuxOut[5] = fifoOut[23][4][w-1];
              unloadMuxOut[6] = fifoOut[24][4][w-1];
              unloadMuxOut[7] = fifoOut[25][4][w-1];
              unloadMuxOut[8] = fifoOut[0][3][w-1];
              unloadMuxOut[9] = fifoOut[1][3][w-1];
              unloadMuxOut[10] = fifoOut[2][3][w-1];
              unloadMuxOut[11] = fifoOut[3][3][w-1];
              unloadMuxOut[12] = fifoOut[4][3][w-1];
              unloadMuxOut[13] = fifoOut[5][3][w-1];
              unloadMuxOut[14] = fifoOut[6][3][w-1];
              unloadMuxOut[15] = fifoOut[7][3][w-1];
              unloadMuxOut[16] = fifoOut[8][3][w-1];
              unloadMuxOut[17] = fifoOut[9][3][w-1];
              unloadMuxOut[18] = fifoOut[10][3][w-1];
              unloadMuxOut[19] = fifoOut[11][3][w-1];
              unloadMuxOut[20] = fifoOut[12][3][w-1];
              unloadMuxOut[21] = fifoOut[13][3][w-1];
              unloadMuxOut[22] = fifoOut[14][3][w-1];
              unloadMuxOut[23] = fifoOut[15][3][w-1];
              unloadMuxOut[24] = fifoOut[16][3][w-1];
              unloadMuxOut[25] = fifoOut[17][3][w-1];
              unloadMuxOut[26] = fifoOut[18][3][w-1];
              unloadMuxOut[27] = fifoOut[19][3][w-1];
              unloadMuxOut[28] = fifoOut[20][3][w-1];
              unloadMuxOut[29] = fifoOut[21][3][w-1];
              unloadMuxOut[30] = fifoOut[22][3][w-1];
              unloadMuxOut[31] = fifoOut[23][3][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[24][4][w-1];
              unloadMuxOut[1] = fifoOut[25][4][w-1];
              unloadMuxOut[2] = fifoOut[0][3][w-1];
              unloadMuxOut[3] = fifoOut[1][3][w-1];
              unloadMuxOut[4] = fifoOut[2][3][w-1];
              unloadMuxOut[5] = fifoOut[3][3][w-1];
              unloadMuxOut[6] = fifoOut[4][3][w-1];
              unloadMuxOut[7] = fifoOut[5][3][w-1];
              unloadMuxOut[8] = fifoOut[6][3][w-1];
              unloadMuxOut[9] = fifoOut[7][3][w-1];
              unloadMuxOut[10] = fifoOut[8][3][w-1];
              unloadMuxOut[11] = fifoOut[9][3][w-1];
              unloadMuxOut[12] = fifoOut[10][3][w-1];
              unloadMuxOut[13] = fifoOut[11][3][w-1];
              unloadMuxOut[14] = fifoOut[12][3][w-1];
              unloadMuxOut[15] = fifoOut[13][3][w-1];
              unloadMuxOut[16] = fifoOut[14][3][w-1];
              unloadMuxOut[17] = fifoOut[15][3][w-1];
              unloadMuxOut[18] = fifoOut[16][3][w-1];
              unloadMuxOut[19] = fifoOut[17][3][w-1];
              unloadMuxOut[20] = fifoOut[18][3][w-1];
              unloadMuxOut[21] = fifoOut[19][3][w-1];
              unloadMuxOut[22] = fifoOut[20][3][w-1];
              unloadMuxOut[23] = fifoOut[21][3][w-1];
              unloadMuxOut[24] = fifoOut[22][3][w-1];
              unloadMuxOut[25] = fifoOut[23][3][w-1];
              unloadMuxOut[26] = fifoOut[24][3][w-1];
              unloadMuxOut[27] = fifoOut[25][3][w-1];
              unloadMuxOut[28] = fifoOut[0][2][w-1];
              unloadMuxOut[29] = fifoOut[1][2][w-1];
              unloadMuxOut[30] = fifoOut[2][2][w-1];
              unloadMuxOut[31] = fifoOut[3][2][w-1];
       end
       16: begin
              unloadMuxOut[0] = fifoOut[4][3][w-1];
              unloadMuxOut[1] = fifoOut[5][3][w-1];
              unloadMuxOut[2] = fifoOut[6][3][w-1];
              unloadMuxOut[3] = fifoOut[7][3][w-1];
              unloadMuxOut[4] = fifoOut[8][3][w-1];
              unloadMuxOut[5] = fifoOut[9][3][w-1];
              unloadMuxOut[6] = fifoOut[10][3][w-1];
              unloadMuxOut[7] = fifoOut[11][3][w-1];
              unloadMuxOut[8] = fifoOut[12][3][w-1];
              unloadMuxOut[9] = fifoOut[13][3][w-1];
              unloadMuxOut[10] = fifoOut[14][3][w-1];
              unloadMuxOut[11] = fifoOut[15][3][w-1];
              unloadMuxOut[12] = fifoOut[16][3][w-1];
              unloadMuxOut[13] = fifoOut[17][3][w-1];
              unloadMuxOut[14] = fifoOut[18][3][w-1];
              unloadMuxOut[15] = fifoOut[19][3][w-1];
              unloadMuxOut[16] = fifoOut[20][3][w-1];
              unloadMuxOut[17] = fifoOut[21][3][w-1];
              unloadMuxOut[18] = fifoOut[22][3][w-1];
              unloadMuxOut[19] = fifoOut[23][3][w-1];
              unloadMuxOut[20] = fifoOut[24][3][w-1];
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0; 
             end
       end
    endcase //unload case end
    case(iteration_0_indicator)
       0: begin
         case(rd_address_case)
         0: begin
              muxOutConnector[0] = fifoOut[25][4];
              muxOutConnector[1] = fifoOut[0][3];
              muxOutConnector[2] = fifoOut[1][3];
              muxOutConnector[3] = fifoOut[2][3];
              muxOutConnector[4] = fifoOut[3][3];
              muxOutConnector[5] = fifoOut[4][3];
              muxOutConnector[6] = fifoOut[5][3];
              muxOutConnector[7] = fifoOut[6][3];
              muxOutConnector[8] = fifoOut[7][3];
              muxOutConnector[9] = fifoOut[8][3];
              muxOutConnector[10] = fifoOut[9][3];
              muxOutConnector[11] = fifoOut[10][3];
              muxOutConnector[12] = fifoOut[11][3];
              muxOutConnector[13] = fifoOut[12][3];
              muxOutConnector[14] = fifoOut[13][3];
              muxOutConnector[15] = fifoOut[14][3];
              muxOutConnector[16] = fifoOut[15][3];
              muxOutConnector[17] = fifoOut[16][3];
              muxOutConnector[18] = fifoOut[17][3];
              muxOutConnector[19] = fifoOut[18][3];
              muxOutConnector[20] = fifoOut[19][3];
              muxOutConnector[21] = fifoOut[20][3];
              muxOutConnector[22] = fifoOut[21][3];
              muxOutConnector[23] = fifoOut[22][3];
              muxOutConnector[24] = fifoOut[23][3];
              muxOutConnector[25] = fifoOut[24][3];
              muxOutConnector[26] = fifoOut[27][6];
              muxOutConnector[27] = fifoOut[28][6];
              muxOutConnector[28] = fifoOut[29][6];
              muxOutConnector[29] = fifoOut[30][6];
              muxOutConnector[30] = fifoOut[31][6];
              muxOutConnector[31] = fifoOut[32][6];
              muxOutConnector[32] = fifoOut[33][6];
              muxOutConnector[33] = fifoOut[34][6];
              muxOutConnector[34] = fifoOut[35][6];
              muxOutConnector[35] = fifoOut[36][6];
              muxOutConnector[36] = fifoOut[37][6];
              muxOutConnector[37] = fifoOut[38][6];
              muxOutConnector[38] = fifoOut[39][6];
              muxOutConnector[39] = fifoOut[40][6];
              muxOutConnector[40] = fifoOut[41][6];
              muxOutConnector[41] = fifoOut[42][6];
              muxOutConnector[42] = fifoOut[43][6];
              muxOutConnector[43] = fifoOut[44][6];
              muxOutConnector[44] = fifoOut[45][6];
              muxOutConnector[45] = fifoOut[46][6];
              muxOutConnector[46] = fifoOut[47][6];
              muxOutConnector[47] = fifoOut[48][6];
              muxOutConnector[48] = fifoOut[49][6];
              muxOutConnector[49] = fifoOut[50][6];
              muxOutConnector[50] = fifoOut[51][6];
              muxOutConnector[51] = fifoOut[26][5];
         end
         1: begin
              muxOutConnector[0] = fifoOut[25][4];
              muxOutConnector[1] = fifoOut[0][3];
              muxOutConnector[2] = fifoOut[1][3];
              muxOutConnector[3] = fifoOut[2][3];
              muxOutConnector[4] = fifoOut[3][3];
              muxOutConnector[5] = fifoOut[4][3];
              muxOutConnector[6] = fifoOut[5][3];
              muxOutConnector[7] = fifoOut[6][3];
              muxOutConnector[8] = fifoOut[7][3];
              muxOutConnector[9] = fifoOut[8][3];
              muxOutConnector[10] = fifoOut[9][3];
              muxOutConnector[11] = fifoOut[10][3];
              muxOutConnector[12] = fifoOut[11][3];
              muxOutConnector[13] = fifoOut[12][3];
              muxOutConnector[14] = fifoOut[13][3];
              muxOutConnector[15] = fifoOut[14][3];
              muxOutConnector[16] = fifoOut[15][3];
              muxOutConnector[17] = fifoOut[16][3];
              muxOutConnector[18] = fifoOut[17][3];
              muxOutConnector[19] = fifoOut[18][3];
              muxOutConnector[20] = fifoOut[19][3];
              muxOutConnector[21] = fifoOut[20][3];
              muxOutConnector[22] = fifoOut[21][3];
              muxOutConnector[23] = fifoOut[22][3];
              muxOutConnector[24] = fifoOut[23][3];
              muxOutConnector[25] = fifoOut[24][3];
              muxOutConnector[26] = fifoOut[27][6];
              muxOutConnector[27] = fifoOut[28][6];
              muxOutConnector[28] = fifoOut[29][6];
              muxOutConnector[29] = fifoOut[30][6];
              muxOutConnector[30] = fifoOut[31][6];
              muxOutConnector[31] = fifoOut[32][6];
              muxOutConnector[32] = fifoOut[33][6];
              muxOutConnector[33] = fifoOut[34][6];
              muxOutConnector[34] = fifoOut[35][6];
              muxOutConnector[35] = fifoOut[36][6];
              muxOutConnector[36] = fifoOut[37][6];
              muxOutConnector[37] = fifoOut[38][6];
              muxOutConnector[38] = fifoOut[39][6];
              muxOutConnector[39] = fifoOut[40][6];
              muxOutConnector[40] = fifoOut[41][6];
              muxOutConnector[41] = fifoOut[42][6];
              muxOutConnector[42] = fifoOut[43][6];
              muxOutConnector[43] = fifoOut[44][6];
              muxOutConnector[44] = fifoOut[45][6];
              muxOutConnector[45] = fifoOut[46][6];
              muxOutConnector[46] = fifoOut[47][6];
              muxOutConnector[47] = fifoOut[48][6];
              muxOutConnector[48] = fifoOut[49][6];
              muxOutConnector[49] = fifoOut[50][6];
              muxOutConnector[50] = fifoOut[51][6];
              muxOutConnector[51] = fifoOut[26][5];
         end
         2: begin
              muxOutConnector[0] = fifoOut[25][4];
              muxOutConnector[1] = fifoOut[0][3];
              muxOutConnector[2] = fifoOut[1][3];
              muxOutConnector[3] = fifoOut[2][3];
              muxOutConnector[4] = fifoOut[3][3];
              muxOutConnector[5] = fifoOut[4][3];
              muxOutConnector[6] = fifoOut[5][3];
              muxOutConnector[7] = fifoOut[6][3];
              muxOutConnector[8] = fifoOut[7][3];
              muxOutConnector[9] = fifoOut[8][3];
              muxOutConnector[10] = fifoOut[9][3];
              muxOutConnector[11] = fifoOut[10][3];
              muxOutConnector[12] = fifoOut[11][3];
              muxOutConnector[13] = fifoOut[12][3];
              muxOutConnector[14] = fifoOut[13][3];
              muxOutConnector[15] = fifoOut[14][3];
              muxOutConnector[16] = fifoOut[15][3];
              muxOutConnector[17] = fifoOut[16][3];
              muxOutConnector[18] = fifoOut[17][3];
              muxOutConnector[19] = fifoOut[18][3];
              muxOutConnector[20] = fifoOut[19][3];
              muxOutConnector[21] = fifoOut[20][3];
              muxOutConnector[22] = fifoOut[21][3];
              muxOutConnector[23] = fifoOut[22][3];
              muxOutConnector[24] = fifoOut[26][13];
              muxOutConnector[25] = fifoOut[27][13];
              muxOutConnector[26] = fifoOut[27][6];
              muxOutConnector[27] = fifoOut[28][6];
              muxOutConnector[28] = fifoOut[29][6];
              muxOutConnector[29] = fifoOut[30][6];
              muxOutConnector[30] = fifoOut[31][6];
              muxOutConnector[31] = fifoOut[32][6];
              muxOutConnector[32] = fifoOut[33][6];
              muxOutConnector[33] = fifoOut[34][6];
              muxOutConnector[34] = fifoOut[35][6];
              muxOutConnector[35] = fifoOut[36][6];
              muxOutConnector[36] = fifoOut[37][6];
              muxOutConnector[37] = fifoOut[38][6];
              muxOutConnector[38] = fifoOut[39][6];
              muxOutConnector[39] = fifoOut[40][6];
              muxOutConnector[40] = fifoOut[41][6];
              muxOutConnector[41] = fifoOut[42][6];
              muxOutConnector[42] = fifoOut[43][6];
              muxOutConnector[43] = fifoOut[44][6];
              muxOutConnector[44] = fifoOut[45][6];
              muxOutConnector[45] = fifoOut[46][6];
              muxOutConnector[46] = fifoOut[47][6];
              muxOutConnector[47] = fifoOut[48][6];
              muxOutConnector[48] = fifoOut[49][6];
              muxOutConnector[49] = fifoOut[50][6];
              muxOutConnector[50] = fifoOut[51][6];
              muxOutConnector[51] = fifoOut[26][5];
         end
         3: begin
              muxOutConnector[0] = fifoOut[28][14];
              muxOutConnector[1] = fifoOut[29][14];
              muxOutConnector[2] = fifoOut[30][14];
              muxOutConnector[3] = fifoOut[31][14];
              muxOutConnector[4] = fifoOut[32][14];
              muxOutConnector[5] = fifoOut[33][14];
              muxOutConnector[6] = fifoOut[34][14];
              muxOutConnector[7] = fifoOut[35][14];
              muxOutConnector[8] = fifoOut[36][14];
              muxOutConnector[9] = fifoOut[37][14];
              muxOutConnector[10] = fifoOut[38][14];
              muxOutConnector[11] = fifoOut[39][14];
              muxOutConnector[12] = fifoOut[40][14];
              muxOutConnector[13] = fifoOut[41][14];
              muxOutConnector[14] = fifoOut[42][14];
              muxOutConnector[15] = fifoOut[43][14];
              muxOutConnector[16] = fifoOut[44][14];
              muxOutConnector[17] = fifoOut[45][14];
              muxOutConnector[18] = fifoOut[46][14];
              muxOutConnector[19] = fifoOut[47][14];
              muxOutConnector[20] = fifoOut[48][14];
              muxOutConnector[21] = fifoOut[49][14];
              muxOutConnector[22] = fifoOut[50][14];
              muxOutConnector[23] = fifoOut[51][14];
              muxOutConnector[24] = fifoOut[26][13];
              muxOutConnector[25] = fifoOut[27][13];
              muxOutConnector[26] = fifoOut[27][6];
              muxOutConnector[27] = fifoOut[28][6];
              muxOutConnector[28] = fifoOut[29][6];
              muxOutConnector[29] = fifoOut[30][6];
              muxOutConnector[30] = fifoOut[31][6];
              muxOutConnector[31] = fifoOut[32][6];
              muxOutConnector[32] = fifoOut[33][6];
              muxOutConnector[33] = fifoOut[34][6];
              muxOutConnector[34] = fifoOut[35][6];
              muxOutConnector[35] = fifoOut[36][6];
              muxOutConnector[36] = fifoOut[37][6];
              muxOutConnector[37] = fifoOut[38][6];
              muxOutConnector[38] = fifoOut[39][6];
              muxOutConnector[39] = fifoOut[40][6];
              muxOutConnector[40] = fifoOut[41][6];
              muxOutConnector[41] = fifoOut[42][6];
              muxOutConnector[42] = fifoOut[43][6];
              muxOutConnector[43] = fifoOut[44][6];
              muxOutConnector[44] = fifoOut[45][6];
              muxOutConnector[45] = fifoOut[0][14];
              muxOutConnector[46] = fifoOut[1][14];
              muxOutConnector[47] = fifoOut[2][14];
              muxOutConnector[48] = fifoOut[3][14];
              muxOutConnector[49] = fifoOut[4][14];
              muxOutConnector[50] = fifoOut[5][14];
              muxOutConnector[51] = fifoOut[6][14];
         end
         4: begin
              muxOutConnector[0] = fifoOut[28][14];
              muxOutConnector[1] = fifoOut[29][14];
              muxOutConnector[2] = fifoOut[30][14];
              muxOutConnector[3] = fifoOut[31][14];
              muxOutConnector[4] = fifoOut[32][14];
              muxOutConnector[5] = fifoOut[33][14];
              muxOutConnector[6] = fifoOut[34][14];
              muxOutConnector[7] = fifoOut[35][14];
              muxOutConnector[8] = fifoOut[36][14];
              muxOutConnector[9] = fifoOut[37][14];
              muxOutConnector[10] = fifoOut[38][14];
              muxOutConnector[11] = fifoOut[39][14];
              muxOutConnector[12] = fifoOut[40][14];
              muxOutConnector[13] = fifoOut[41][14];
              muxOutConnector[14] = fifoOut[42][14];
              muxOutConnector[15] = fifoOut[43][14];
              muxOutConnector[16] = fifoOut[44][14];
              muxOutConnector[17] = fifoOut[45][14];
              muxOutConnector[18] = fifoOut[46][14];
              muxOutConnector[19] = fifoOut[47][14];
              muxOutConnector[20] = fifoOut[48][14];
              muxOutConnector[21] = fifoOut[49][14];
              muxOutConnector[22] = fifoOut[50][14];
              muxOutConnector[23] = fifoOut[51][14];
              muxOutConnector[24] = fifoOut[26][13];
              muxOutConnector[25] = fifoOut[27][13];
              muxOutConnector[26] = fifoOut[7][15];
              muxOutConnector[27] = fifoOut[8][15];
              muxOutConnector[28] = fifoOut[9][15];
              muxOutConnector[29] = fifoOut[10][15];
              muxOutConnector[30] = fifoOut[11][15];
              muxOutConnector[31] = fifoOut[12][15];
              muxOutConnector[32] = fifoOut[13][15];
              muxOutConnector[33] = fifoOut[14][15];
              muxOutConnector[34] = fifoOut[15][15];
              muxOutConnector[35] = fifoOut[16][15];
              muxOutConnector[36] = fifoOut[17][15];
              muxOutConnector[37] = fifoOut[18][15];
              muxOutConnector[38] = fifoOut[19][15];
              muxOutConnector[39] = fifoOut[20][15];
              muxOutConnector[40] = fifoOut[21][15];
              muxOutConnector[41] = fifoOut[22][15];
              muxOutConnector[42] = fifoOut[23][15];
              muxOutConnector[43] = fifoOut[24][15];
              muxOutConnector[44] = fifoOut[25][15];
              muxOutConnector[45] = fifoOut[0][14];
              muxOutConnector[46] = fifoOut[1][14];
              muxOutConnector[47] = fifoOut[2][14];
              muxOutConnector[48] = fifoOut[3][14];
              muxOutConnector[49] = fifoOut[4][14];
              muxOutConnector[50] = fifoOut[5][14];
              muxOutConnector[51] = fifoOut[6][14];
         end
         5: begin
              muxOutConnector[0] = fifoOut[28][14];
              muxOutConnector[1] = fifoOut[29][14];
              muxOutConnector[2] = fifoOut[30][14];
              muxOutConnector[3] = fifoOut[31][14];
              muxOutConnector[4] = fifoOut[32][14];
              muxOutConnector[5] = fifoOut[33][14];
              muxOutConnector[6] = fifoOut[34][14];
              muxOutConnector[7] = fifoOut[35][14];
              muxOutConnector[8] = fifoOut[36][14];
              muxOutConnector[9] = fifoOut[37][14];
              muxOutConnector[10] = fifoOut[38][14];
              muxOutConnector[11] = fifoOut[39][14];
              muxOutConnector[12] = fifoOut[40][14];
              muxOutConnector[13] = fifoOut[41][14];
              muxOutConnector[14] = fifoOut[42][14];
              muxOutConnector[15] = fifoOut[43][14];
              muxOutConnector[16] = fifoOut[44][14];
              muxOutConnector[17] = fifoOut[45][14];
              muxOutConnector[18] = fifoOut[46][14];
              muxOutConnector[19] = fifoOut[47][14];
              muxOutConnector[20] = fifoOut[48][14];
              muxOutConnector[21] = fifoOut[49][14];
              muxOutConnector[22] = fifoOut[50][14];
              muxOutConnector[23] = fifoOut[51][14];
              muxOutConnector[24] = fifoOut[26][13];
              muxOutConnector[25] = fifoOut[27][13];
              muxOutConnector[26] = fifoOut[7][15];
              muxOutConnector[27] = fifoOut[8][15];
              muxOutConnector[28] = fifoOut[9][15];
              muxOutConnector[29] = fifoOut[10][15];
              muxOutConnector[30] = fifoOut[11][15];
              muxOutConnector[31] = fifoOut[12][15];
              muxOutConnector[32] = fifoOut[13][15];
              muxOutConnector[33] = fifoOut[14][15];
              muxOutConnector[34] = fifoOut[15][15];
              muxOutConnector[35] = fifoOut[16][15];
              muxOutConnector[36] = fifoOut[17][15];
              muxOutConnector[37] = fifoOut[18][15];
              muxOutConnector[38] = fifoOut[19][15];
              muxOutConnector[39] = fifoOut[20][15];
              muxOutConnector[40] = fifoOut[21][15];
              muxOutConnector[41] = fifoOut[22][15];
              muxOutConnector[42] = fifoOut[23][15];
              muxOutConnector[43] = fifoOut[24][15];
              muxOutConnector[44] = fifoOut[25][15];
              muxOutConnector[45] = fifoOut[0][14];
              muxOutConnector[46] = fifoOut[1][14];
              muxOutConnector[47] = fifoOut[2][14];
              muxOutConnector[48] = fifoOut[3][14];
              muxOutConnector[49] = fifoOut[4][14];
              muxOutConnector[50] = fifoOut[5][14];
              muxOutConnector[51] = fifoOut[6][14];
         end
         6: begin
              muxOutConnector[0] = fifoOut[28][14];
              muxOutConnector[1] = fifoOut[29][14];
              muxOutConnector[2] = fifoOut[30][14];
              muxOutConnector[3] = fifoOut[31][14];
              muxOutConnector[4] = fifoOut[32][14];
              muxOutConnector[5] = fifoOut[33][14];
              muxOutConnector[6] = fifoOut[34][14];
              muxOutConnector[7] = fifoOut[35][14];
              muxOutConnector[8] = fifoOut[36][14];
              muxOutConnector[9] = fifoOut[37][14];
              muxOutConnector[10] = fifoOut[38][14];
              muxOutConnector[11] = fifoOut[39][14];
              muxOutConnector[12] = fifoOut[40][14];
              muxOutConnector[13] = fifoOut[41][14];
              muxOutConnector[14] = fifoOut[42][14];
              muxOutConnector[15] = fifoOut[43][14];
              muxOutConnector[16] = fifoOut[44][14];
              muxOutConnector[17] = fifoOut[45][14];
              muxOutConnector[18] = fifoOut[46][14];
              muxOutConnector[19] = fifoOut[47][14];
              muxOutConnector[20] = fifoOut[48][14];
              muxOutConnector[21] = fifoOut[49][14];
              muxOutConnector[22] = fifoOut[50][14];
              muxOutConnector[23] = fifoOut[51][14];
              muxOutConnector[24] = fifoOut[26][13];
              muxOutConnector[25] = fifoOut[27][13];
              muxOutConnector[26] = fifoOut[7][15];
              muxOutConnector[27] = fifoOut[8][15];
              muxOutConnector[28] = fifoOut[9][15];
              muxOutConnector[29] = fifoOut[10][15];
              muxOutConnector[30] = fifoOut[11][15];
              muxOutConnector[31] = fifoOut[12][15];
              muxOutConnector[32] = fifoOut[13][15];
              muxOutConnector[33] = fifoOut[14][15];
              muxOutConnector[34] = fifoOut[15][15];
              muxOutConnector[35] = fifoOut[16][15];
              muxOutConnector[36] = fifoOut[17][15];
              muxOutConnector[37] = fifoOut[18][15];
              muxOutConnector[38] = fifoOut[19][15];
              muxOutConnector[39] = fifoOut[20][15];
              muxOutConnector[40] = fifoOut[21][15];
              muxOutConnector[41] = fifoOut[22][15];
              muxOutConnector[42] = fifoOut[23][15];
              muxOutConnector[43] = fifoOut[24][15];
              muxOutConnector[44] = fifoOut[25][15];
              muxOutConnector[45] = fifoOut[0][14];
              muxOutConnector[46] = fifoOut[1][14];
              muxOutConnector[47] = fifoOut[2][14];
              muxOutConnector[48] = fifoOut[3][14];
              muxOutConnector[49] = fifoOut[4][14];
              muxOutConnector[50] = fifoOut[5][14];
              muxOutConnector[51] = fifoOut[6][14];
         end
         7: begin
              muxOutConnector[0] = fifoOut[28][14];
              muxOutConnector[1] = fifoOut[29][14];
              muxOutConnector[2] = fifoOut[30][14];
              muxOutConnector[3] = fifoOut[31][14];
              muxOutConnector[4] = fifoOut[32][14];
              muxOutConnector[5] = fifoOut[33][14];
              muxOutConnector[6] = fifoOut[34][14];
              muxOutConnector[7] = fifoOut[35][14];
              muxOutConnector[8] = fifoOut[36][14];
              muxOutConnector[9] = fifoOut[37][14];
              muxOutConnector[10] = fifoOut[38][14];
              muxOutConnector[11] = fifoOut[39][14];
              muxOutConnector[12] = fifoOut[40][14];
              muxOutConnector[13] = fifoOut[41][14];
              muxOutConnector[14] = fifoOut[42][14];
              muxOutConnector[15] = fifoOut[43][14];
              muxOutConnector[16] = fifoOut[44][14];
              muxOutConnector[17] = fifoOut[45][14];
              muxOutConnector[18] = fifoOut[46][14];
              muxOutConnector[19] = fifoOut[47][14];
              muxOutConnector[20] = fifoOut[48][14];
              muxOutConnector[21] = fifoOut[49][14];
              muxOutConnector[22] = fifoOut[50][14];
              muxOutConnector[23] = fifoOut[51][14];
              muxOutConnector[24] = fifoOut[26][13];
              muxOutConnector[25] = fifoOut[27][13];
              muxOutConnector[26] = fifoOut[7][15];
              muxOutConnector[27] = fifoOut[8][15];
              muxOutConnector[28] = fifoOut[9][15];
              muxOutConnector[29] = fifoOut[10][15];
              muxOutConnector[30] = fifoOut[11][15];
              muxOutConnector[31] = fifoOut[12][15];
              muxOutConnector[32] = fifoOut[13][15];
              muxOutConnector[33] = fifoOut[14][15];
              muxOutConnector[34] = fifoOut[15][15];
              muxOutConnector[35] = fifoOut[16][15];
              muxOutConnector[36] = fifoOut[17][15];
              muxOutConnector[37] = fifoOut[18][15];
              muxOutConnector[38] = fifoOut[19][15];
              muxOutConnector[39] = fifoOut[20][15];
              muxOutConnector[40] = fifoOut[21][15];
              muxOutConnector[41] = fifoOut[22][15];
              muxOutConnector[42] = fifoOut[23][15];
              muxOutConnector[43] = fifoOut[24][15];
              muxOutConnector[44] = fifoOut[25][15];
              muxOutConnector[45] = fifoOut[0][14];
              muxOutConnector[46] = fifoOut[1][14];
              muxOutConnector[47] = fifoOut[2][14];
              muxOutConnector[48] = fifoOut[3][14];
              muxOutConnector[49] = fifoOut[4][14];
              muxOutConnector[50] = fifoOut[5][14];
              muxOutConnector[51] = fifoOut[6][14];
         end
         8: begin
              muxOutConnector[0] = fifoOut[28][14];
              muxOutConnector[1] = fifoOut[29][14];
              muxOutConnector[2] = fifoOut[30][14];
              muxOutConnector[3] = fifoOut[31][14];
              muxOutConnector[4] = fifoOut[32][14];
              muxOutConnector[5] = fifoOut[33][14];
              muxOutConnector[6] = fifoOut[34][14];
              muxOutConnector[7] = fifoOut[35][14];
              muxOutConnector[8] = fifoOut[36][14];
              muxOutConnector[9] = fifoOut[37][14];
              muxOutConnector[10] = fifoOut[38][14];
              muxOutConnector[11] = fifoOut[39][14];
              muxOutConnector[12] = fifoOut[40][14];
              muxOutConnector[13] = fifoOut[41][14];
              muxOutConnector[14] = fifoOut[42][14];
              muxOutConnector[15] = fifoOut[43][14];
              muxOutConnector[16] = fifoOut[44][14];
              muxOutConnector[17] = fifoOut[45][14];
              muxOutConnector[18] = fifoOut[46][14];
              muxOutConnector[19] = fifoOut[47][14];
              muxOutConnector[20] = fifoOut[48][14];
              muxOutConnector[21] = fifoOut[49][14];
              muxOutConnector[22] = fifoOut[50][14];
              muxOutConnector[23] = fifoOut[51][14];
              muxOutConnector[24] = fifoOut[26][13];
              muxOutConnector[25] = fifoOut[27][13];
              muxOutConnector[26] = fifoOut[7][15];
              muxOutConnector[27] = fifoOut[8][15];
              muxOutConnector[28] = fifoOut[9][15];
              muxOutConnector[29] = fifoOut[10][15];
              muxOutConnector[30] = fifoOut[11][15];
              muxOutConnector[31] = fifoOut[12][15];
              muxOutConnector[32] = fifoOut[13][15];
              muxOutConnector[33] = fifoOut[14][15];
              muxOutConnector[34] = fifoOut[15][15];
              muxOutConnector[35] = fifoOut[16][15];
              muxOutConnector[36] = fifoOut[17][15];
              muxOutConnector[37] = fifoOut[18][15];
              muxOutConnector[38] = fifoOut[19][15];
              muxOutConnector[39] = fifoOut[20][15];
              muxOutConnector[40] = fifoOut[21][15];
              muxOutConnector[41] = fifoOut[22][15];
              muxOutConnector[42] = fifoOut[23][15];
              muxOutConnector[43] = fifoOut[24][15];
              muxOutConnector[44] = fifoOut[25][15];
              muxOutConnector[45] = fifoOut[0][14];
              muxOutConnector[46] = fifoOut[1][14];
              muxOutConnector[47] = fifoOut[2][14];
              muxOutConnector[48] = fifoOut[3][14];
              muxOutConnector[49] = fifoOut[4][14];
              muxOutConnector[50] = fifoOut[5][14];
              muxOutConnector[51] = fifoOut[6][14];
         end
         9: begin
              muxOutConnector[0] = fifoOut[28][14];
              muxOutConnector[1] = fifoOut[29][14];
              muxOutConnector[2] = fifoOut[30][14];
              muxOutConnector[3] = fifoOut[31][14];
              muxOutConnector[4] = fifoOut[32][14];
              muxOutConnector[5] = fifoOut[33][14];
              muxOutConnector[6] = fifoOut[34][14];
              muxOutConnector[7] = fifoOut[35][14];
              muxOutConnector[8] = fifoOut[36][14];
              muxOutConnector[9] = fifoOut[37][14];
              muxOutConnector[10] = fifoOut[38][14];
              muxOutConnector[11] = fifoOut[39][14];
              muxOutConnector[12] = fifoOut[40][14];
              muxOutConnector[13] = fifoOut[41][14];
              muxOutConnector[14] = fifoOut[42][14];
              muxOutConnector[15] = fifoOut[43][14];
              muxOutConnector[16] = fifoOut[44][14];
              muxOutConnector[17] = fifoOut[45][14];
              muxOutConnector[18] = fifoOut[46][14];
              muxOutConnector[19] = fifoOut[47][14];
              muxOutConnector[20] = fifoOut[48][14];
              muxOutConnector[21] = fifoOut[49][14];
              muxOutConnector[22] = fifoOut[50][14];
              muxOutConnector[23] = fifoOut[51][14];
              muxOutConnector[24] = fifoOut[26][13];
              muxOutConnector[25] = fifoOut[27][13];
              muxOutConnector[26] = fifoOut[7][15];
              muxOutConnector[27] = fifoOut[8][15];
              muxOutConnector[28] = fifoOut[9][15];
              muxOutConnector[29] = fifoOut[10][15];
              muxOutConnector[30] = fifoOut[11][15];
              muxOutConnector[31] = fifoOut[12][15];
              muxOutConnector[32] = fifoOut[13][15];
              muxOutConnector[33] = fifoOut[14][15];
              muxOutConnector[34] = fifoOut[15][15];
              muxOutConnector[35] = fifoOut[16][15];
              muxOutConnector[36] = fifoOut[17][15];
              muxOutConnector[37] = fifoOut[18][15];
              muxOutConnector[38] = fifoOut[19][15];
              muxOutConnector[39] = fifoOut[20][15];
              muxOutConnector[40] = fifoOut[21][15];
              muxOutConnector[41] = fifoOut[22][15];
              muxOutConnector[42] = fifoOut[23][15];
              muxOutConnector[43] = fifoOut[24][15];
              muxOutConnector[44] = fifoOut[25][15];
              muxOutConnector[45] = fifoOut[0][14];
              muxOutConnector[46] = fifoOut[1][14];
              muxOutConnector[47] = fifoOut[2][14];
              muxOutConnector[48] = fifoOut[3][14];
              muxOutConnector[49] = fifoOut[4][14];
              muxOutConnector[50] = fifoOut[5][14];
              muxOutConnector[51] = fifoOut[6][14];
         end
         10: begin
              muxOutConnector[0] = fifoOut[28][14];
              muxOutConnector[1] = fifoOut[29][14];
              muxOutConnector[2] = fifoOut[30][14];
              muxOutConnector[3] = fifoOut[31][14];
              muxOutConnector[4] = fifoOut[32][14];
              muxOutConnector[5] = fifoOut[33][14];
              muxOutConnector[6] = fifoOut[34][14];
              muxOutConnector[7] = fifoOut[35][14];
              muxOutConnector[8] = fifoOut[36][14];
              muxOutConnector[9] = fifoOut[37][14];
              muxOutConnector[10] = fifoOut[38][14];
              muxOutConnector[11] = fifoOut[39][14];
              muxOutConnector[12] = fifoOut[40][14];
              muxOutConnector[13] = fifoOut[41][14];
              muxOutConnector[14] = fifoOut[42][14];
              muxOutConnector[15] = fifoOut[43][14];
              muxOutConnector[16] = fifoOut[44][14];
              muxOutConnector[17] = fifoOut[45][14];
              muxOutConnector[18] = fifoOut[46][14];
              muxOutConnector[19] = fifoOut[47][14];
              muxOutConnector[20] = fifoOut[48][14];
              muxOutConnector[21] = fifoOut[49][14];
              muxOutConnector[22] = fifoOut[50][14];
              muxOutConnector[23] = fifoOut[51][14];
              muxOutConnector[24] = fifoOut[26][13];
              muxOutConnector[25] = fifoOut[27][13];
              muxOutConnector[26] = fifoOut[7][15];
              muxOutConnector[27] = fifoOut[8][15];
              muxOutConnector[28] = fifoOut[9][15];
              muxOutConnector[29] = fifoOut[10][15];
              muxOutConnector[30] = fifoOut[11][15];
              muxOutConnector[31] = fifoOut[12][15];
              muxOutConnector[32] = fifoOut[13][15];
              muxOutConnector[33] = fifoOut[14][15];
              muxOutConnector[34] = fifoOut[15][15];
              muxOutConnector[35] = fifoOut[16][15];
              muxOutConnector[36] = fifoOut[17][15];
              muxOutConnector[37] = fifoOut[18][15];
              muxOutConnector[38] = fifoOut[19][15];
              muxOutConnector[39] = fifoOut[20][15];
              muxOutConnector[40] = fifoOut[21][15];
              muxOutConnector[41] = fifoOut[22][15];
              muxOutConnector[42] = fifoOut[23][15];
              muxOutConnector[43] = fifoOut[24][15];
              muxOutConnector[44] = fifoOut[25][15];
              muxOutConnector[45] = fifoOut[0][14];
              muxOutConnector[46] = fifoOut[1][14];
              muxOutConnector[47] = fifoOut[2][14];
              muxOutConnector[48] = fifoOut[3][14];
              muxOutConnector[49] = fifoOut[4][14];
              muxOutConnector[50] = fifoOut[5][14];
              muxOutConnector[51] = fifoOut[6][14];
         end
         11: begin
              muxOutConnector[0] = fifoOut[28][14];
              muxOutConnector[1] = fifoOut[29][14];
              muxOutConnector[2] = fifoOut[30][14];
              muxOutConnector[3] = fifoOut[31][14];
              muxOutConnector[4] = fifoOut[32][14];
              muxOutConnector[5] = fifoOut[33][14];
              muxOutConnector[6] = fifoOut[34][14];
              muxOutConnector[7] = fifoOut[35][14];
              muxOutConnector[8] = fifoOut[36][14];
              muxOutConnector[9] = fifoOut[37][14];
              muxOutConnector[10] = fifoOut[38][14];
              muxOutConnector[11] = fifoOut[39][14];
              muxOutConnector[12] = fifoOut[40][14];
              muxOutConnector[13] = fifoOut[41][14];
              muxOutConnector[14] = fifoOut[42][14];
              muxOutConnector[15] = fifoOut[43][14];
              muxOutConnector[16] = fifoOut[44][14];
              muxOutConnector[17] = fifoOut[45][14];
              muxOutConnector[18] = fifoOut[46][14];
              muxOutConnector[19] = fifoOut[47][14];
              muxOutConnector[20] = fifoOut[48][14];
              muxOutConnector[21] = fifoOut[49][14];
              muxOutConnector[22] = fifoOut[50][14];
              muxOutConnector[23] = fifoOut[51][14];
              muxOutConnector[24] = fifoOut[26][13];
              muxOutConnector[25] = fifoOut[27][13];
              muxOutConnector[26] = fifoOut[7][15];
              muxOutConnector[27] = fifoOut[8][15];
              muxOutConnector[28] = fifoOut[9][15];
              muxOutConnector[29] = fifoOut[10][15];
              muxOutConnector[30] = fifoOut[11][15];
              muxOutConnector[31] = fifoOut[12][15];
              muxOutConnector[32] = fifoOut[13][15];
              muxOutConnector[33] = fifoOut[14][15];
              muxOutConnector[34] = fifoOut[15][15];
              muxOutConnector[35] = fifoOut[16][15];
              muxOutConnector[36] = fifoOut[17][15];
              muxOutConnector[37] = fifoOut[18][15];
              muxOutConnector[38] = fifoOut[19][15];
              muxOutConnector[39] = fifoOut[20][15];
              muxOutConnector[40] = fifoOut[21][15];
              muxOutConnector[41] = fifoOut[22][15];
              muxOutConnector[42] = fifoOut[23][15];
              muxOutConnector[43] = fifoOut[24][15];
              muxOutConnector[44] = fifoOut[25][15];
              muxOutConnector[45] = fifoOut[0][14];
              muxOutConnector[46] = fifoOut[1][14];
              muxOutConnector[47] = fifoOut[2][14];
              muxOutConnector[48] = fifoOut[3][14];
              muxOutConnector[49] = fifoOut[4][14];
              muxOutConnector[50] = fifoOut[5][14];
              muxOutConnector[51] = fifoOut[6][14];
         end
         12: begin
              muxOutConnector[0] = fifoOut[28][14];
              muxOutConnector[1] = fifoOut[29][14];
              muxOutConnector[2] = fifoOut[30][14];
              muxOutConnector[3] = fifoOut[31][14];
              muxOutConnector[4] = fifoOut[32][14];
              muxOutConnector[5] = fifoOut[33][14];
              muxOutConnector[6] = fifoOut[34][14];
              muxOutConnector[7] = fifoOut[35][14];
              muxOutConnector[8] = fifoOut[36][14];
              muxOutConnector[9] = fifoOut[37][14];
              muxOutConnector[10] = fifoOut[38][14];
              muxOutConnector[11] = fifoOut[39][14];
              muxOutConnector[12] = fifoOut[40][14];
              muxOutConnector[13] = fifoOut[41][14];
              muxOutConnector[14] = fifoOut[42][14];
              muxOutConnector[15] = fifoOut[43][14];
              muxOutConnector[16] = fifoOut[44][14];
              muxOutConnector[17] = fifoOut[45][14];
              muxOutConnector[18] = fifoOut[46][14];
              muxOutConnector[19] = fifoOut[47][14];
              muxOutConnector[20] = fifoOut[48][14];
              muxOutConnector[21] = fifoOut[49][14];
              muxOutConnector[22] = fifoOut[50][14];
              muxOutConnector[23] = fifoOut[51][14];
              muxOutConnector[24] = fifoOut[26][13];
              muxOutConnector[25] = fifoOut[27][13];
              muxOutConnector[26] = fifoOut[7][15];
              muxOutConnector[27] = fifoOut[8][15];
              muxOutConnector[28] = fifoOut[9][15];
              muxOutConnector[29] = fifoOut[10][15];
              muxOutConnector[30] = fifoOut[11][15];
              muxOutConnector[31] = fifoOut[12][15];
              muxOutConnector[32] = fifoOut[13][15];
              muxOutConnector[33] = fifoOut[14][15];
              muxOutConnector[34] = fifoOut[15][15];
              muxOutConnector[35] = fifoOut[16][15];
              muxOutConnector[36] = fifoOut[17][15];
              muxOutConnector[37] = fifoOut[18][15];
              muxOutConnector[38] = fifoOut[19][15];
              muxOutConnector[39] = fifoOut[20][15];
              muxOutConnector[40] = fifoOut[21][15];
              muxOutConnector[41] = fifoOut[22][15];
              muxOutConnector[42] = fifoOut[23][15];
              muxOutConnector[43] = fifoOut[24][15];
              muxOutConnector[44] = fifoOut[25][15];
              muxOutConnector[45] = fifoOut[0][14];
              muxOutConnector[46] = fifoOut[1][14];
              muxOutConnector[47] = fifoOut[2][14];
              muxOutConnector[48] = fifoOut[3][14];
              muxOutConnector[49] = fifoOut[4][14];
              muxOutConnector[50] = fifoOut[5][14];
              muxOutConnector[51] = fifoOut[6][14];
         end
         13: begin
              muxOutConnector[0] = fifoOut[28][14];
              muxOutConnector[1] = fifoOut[29][14];
              muxOutConnector[2] = fifoOut[30][14];
              muxOutConnector[3] = fifoOut[31][14];
              muxOutConnector[4] = fifoOut[32][14];
              muxOutConnector[5] = fifoOut[33][14];
              muxOutConnector[6] = fifoOut[34][14];
              muxOutConnector[7] = fifoOut[35][14];
              muxOutConnector[8] = fifoOut[36][14];
              muxOutConnector[9] = fifoOut[37][14];
              muxOutConnector[10] = fifoOut[38][14];
              muxOutConnector[11] = fifoOut[39][14];
              muxOutConnector[12] = fifoOut[40][14];
              muxOutConnector[13] = fifoOut[41][14];
              muxOutConnector[14] = fifoOut[42][14];
              muxOutConnector[15] = fifoOut[43][14];
              muxOutConnector[16] = fifoOut[44][14];
              muxOutConnector[17] = fifoOut[45][14];
              muxOutConnector[18] = fifoOut[46][14];
              muxOutConnector[19] = fifoOut[47][14];
              muxOutConnector[20] = fifoOut[48][14];
              muxOutConnector[21] = fifoOut[49][14];
              muxOutConnector[22] = fifoOut[50][14];
              muxOutConnector[23] = fifoOut[51][14];
              muxOutConnector[24] = fifoOut[26][13];
              muxOutConnector[25] = fifoOut[27][13];
              muxOutConnector[26] = fifoOut[7][15];
              muxOutConnector[27] = fifoOut[8][15];
              muxOutConnector[28] = fifoOut[9][15];
              muxOutConnector[29] = fifoOut[10][15];
              muxOutConnector[30] = fifoOut[11][15];
              muxOutConnector[31] = fifoOut[12][15];
              muxOutConnector[32] = fifoOut[13][15];
              muxOutConnector[33] = fifoOut[14][15];
              muxOutConnector[34] = fifoOut[15][15];
              muxOutConnector[35] = fifoOut[16][15];
              muxOutConnector[36] = fifoOut[17][15];
              muxOutConnector[37] = fifoOut[18][15];
              muxOutConnector[38] = fifoOut[19][15];
              muxOutConnector[39] = fifoOut[20][15];
              muxOutConnector[40] = fifoOut[21][15];
              muxOutConnector[41] = fifoOut[22][15];
              muxOutConnector[42] = fifoOut[23][15];
              muxOutConnector[43] = fifoOut[24][15];
              muxOutConnector[44] = fifoOut[25][15];
              muxOutConnector[45] = fifoOut[0][14];
              muxOutConnector[46] = fifoOut[1][14];
              muxOutConnector[47] = fifoOut[2][14];
              muxOutConnector[48] = fifoOut[3][14];
              muxOutConnector[49] = fifoOut[4][14];
              muxOutConnector[50] = fifoOut[5][14];
              muxOutConnector[51] = fifoOut[6][14];
         end
         14: begin
              muxOutConnector[0] = fifoOut[28][14];
              muxOutConnector[1] = fifoOut[29][14];
              muxOutConnector[2] = fifoOut[30][14];
              muxOutConnector[3] = fifoOut[31][14];
              muxOutConnector[4] = fifoOut[32][14];
              muxOutConnector[5] = fifoOut[33][14];
              muxOutConnector[6] = fifoOut[34][14];
              muxOutConnector[7] = fifoOut[35][14];
              muxOutConnector[8] = fifoOut[36][14];
              muxOutConnector[9] = fifoOut[37][14];
              muxOutConnector[10] = fifoOut[38][14];
              muxOutConnector[11] = fifoOut[39][14];
              muxOutConnector[12] = fifoOut[40][14];
              muxOutConnector[13] = fifoOut[41][14];
              muxOutConnector[14] = fifoOut[42][14];
              muxOutConnector[15] = fifoOut[23][6];
              muxOutConnector[16] = fifoOut[24][6];
              muxOutConnector[17] = fifoOut[25][6];
              muxOutConnector[18] = fifoOut[0][5];
              muxOutConnector[19] = fifoOut[1][5];
              muxOutConnector[20] = fifoOut[2][5];
              muxOutConnector[21] = fifoOut[3][5];
              muxOutConnector[22] = fifoOut[4][5];
              muxOutConnector[23] = fifoOut[5][5];
              muxOutConnector[24] = fifoOut[6][5];
              muxOutConnector[25] = fifoOut[7][5];
              muxOutConnector[26] = fifoOut[7][15];
              muxOutConnector[27] = fifoOut[8][15];
              muxOutConnector[28] = fifoOut[9][15];
              muxOutConnector[29] = fifoOut[10][15];
              muxOutConnector[30] = fifoOut[11][15];
              muxOutConnector[31] = fifoOut[12][15];
              muxOutConnector[32] = fifoOut[13][15];
              muxOutConnector[33] = fifoOut[14][15];
              muxOutConnector[34] = fifoOut[15][15];
              muxOutConnector[35] = fifoOut[16][15];
              muxOutConnector[36] = fifoOut[17][15];
              muxOutConnector[37] = fifoOut[18][15];
              muxOutConnector[38] = fifoOut[19][15];
              muxOutConnector[39] = fifoOut[20][15];
              muxOutConnector[40] = fifoOut[21][15];
              muxOutConnector[41] = fifoOut[22][15];
              muxOutConnector[42] = fifoOut[23][15];
              muxOutConnector[43] = fifoOut[24][15];
              muxOutConnector[44] = fifoOut[25][15];
              muxOutConnector[45] = fifoOut[0][14];
              muxOutConnector[46] = fifoOut[1][14];
              muxOutConnector[47] = fifoOut[2][14];
              muxOutConnector[48] = fifoOut[3][14];
              muxOutConnector[49] = fifoOut[4][14];
              muxOutConnector[50] = fifoOut[5][14];
              muxOutConnector[51] = fifoOut[6][14];
         end
         15: begin
              muxOutConnector[0] = fifoOut[8][6];
              muxOutConnector[1] = fifoOut[9][6];
              muxOutConnector[2] = fifoOut[10][6];
              muxOutConnector[3] = fifoOut[11][6];
              muxOutConnector[4] = fifoOut[12][6];
              muxOutConnector[5] = fifoOut[13][6];
              muxOutConnector[6] = fifoOut[14][6];
              muxOutConnector[7] = fifoOut[15][6];
              muxOutConnector[8] = fifoOut[16][6];
              muxOutConnector[9] = fifoOut[17][6];
              muxOutConnector[10] = fifoOut[18][6];
              muxOutConnector[11] = fifoOut[19][6];
              muxOutConnector[12] = fifoOut[20][6];
              muxOutConnector[13] = fifoOut[21][6];
              muxOutConnector[14] = fifoOut[22][6];
              muxOutConnector[15] = fifoOut[23][6];
              muxOutConnector[16] = fifoOut[24][6];
              muxOutConnector[17] = fifoOut[25][6];
              muxOutConnector[18] = fifoOut[0][5];
              muxOutConnector[19] = fifoOut[1][5];
              muxOutConnector[20] = fifoOut[2][5];
              muxOutConnector[21] = fifoOut[3][5];
              muxOutConnector[22] = fifoOut[4][5];
              muxOutConnector[23] = fifoOut[5][5];
              muxOutConnector[24] = fifoOut[6][5];
              muxOutConnector[25] = fifoOut[7][5];
              muxOutConnector[26] = fifoOut[7][15];
              muxOutConnector[27] = fifoOut[8][15];
              muxOutConnector[28] = fifoOut[9][15];
              muxOutConnector[29] = fifoOut[10][15];
              muxOutConnector[30] = fifoOut[11][15];
              muxOutConnector[31] = fifoOut[12][15];
              muxOutConnector[32] = fifoOut[13][15];
              muxOutConnector[33] = fifoOut[14][15];
              muxOutConnector[34] = fifoOut[15][15];
              muxOutConnector[35] = fifoOut[16][15];
              muxOutConnector[36] = fifoOut[46][9];
              muxOutConnector[37] = fifoOut[47][9];
              muxOutConnector[38] = fifoOut[48][9];
              muxOutConnector[39] = fifoOut[49][9];
              muxOutConnector[40] = fifoOut[50][9];
              muxOutConnector[41] = fifoOut[51][9];
              muxOutConnector[42] = fifoOut[26][8];
              muxOutConnector[43] = fifoOut[27][8];
              muxOutConnector[44] = fifoOut[28][8];
              muxOutConnector[45] = fifoOut[29][8];
              muxOutConnector[46] = fifoOut[30][8];
              muxOutConnector[47] = fifoOut[31][8];
              muxOutConnector[48] = fifoOut[32][8];
              muxOutConnector[49] = fifoOut[33][8];
              muxOutConnector[50] = fifoOut[34][8];
              muxOutConnector[51] = fifoOut[35][8];
         end
         16: begin
              muxOutConnector[0] = fifoOut[8][6];
              muxOutConnector[1] = fifoOut[9][6];
              muxOutConnector[2] = fifoOut[10][6];
              muxOutConnector[3] = fifoOut[11][6];
              muxOutConnector[4] = fifoOut[12][6];
              muxOutConnector[5] = fifoOut[13][6];
              muxOutConnector[6] = fifoOut[14][6];
              muxOutConnector[7] = fifoOut[15][6];
              muxOutConnector[8] = fifoOut[16][6];
              muxOutConnector[9] = fifoOut[17][6];
              muxOutConnector[10] = fifoOut[18][6];
              muxOutConnector[11] = fifoOut[19][6];
              muxOutConnector[12] = fifoOut[20][6];
              muxOutConnector[13] = fifoOut[21][6];
              muxOutConnector[14] = fifoOut[22][6];
              muxOutConnector[15] = fifoOut[23][6];
              muxOutConnector[16] = fifoOut[24][6];
              muxOutConnector[17] = fifoOut[25][6];
              muxOutConnector[18] = fifoOut[0][5];
              muxOutConnector[19] = fifoOut[1][5];
              muxOutConnector[20] = fifoOut[2][5];
              muxOutConnector[21] = fifoOut[3][5];
              muxOutConnector[22] = fifoOut[4][5];
              muxOutConnector[23] = fifoOut[5][5];
              muxOutConnector[24] = fifoOut[6][5];
              muxOutConnector[25] = fifoOut[7][5];
              muxOutConnector[26] = fifoOut[36][9];
              muxOutConnector[27] = fifoOut[37][9];
              muxOutConnector[28] = fifoOut[38][9];
              muxOutConnector[29] = fifoOut[39][9];
              muxOutConnector[30] = fifoOut[40][9];
              muxOutConnector[31] = fifoOut[41][9];
              muxOutConnector[32] = fifoOut[42][9];
              muxOutConnector[33] = fifoOut[43][9];
              muxOutConnector[34] = fifoOut[44][9];
              muxOutConnector[35] = fifoOut[45][9];
              muxOutConnector[36] = fifoOut[46][9];
              muxOutConnector[37] = fifoOut[47][9];
              muxOutConnector[38] = fifoOut[48][9];
              muxOutConnector[39] = fifoOut[49][9];
              muxOutConnector[40] = fifoOut[50][9];
              muxOutConnector[41] = fifoOut[51][9];
              muxOutConnector[42] = fifoOut[26][8];
              muxOutConnector[43] = fifoOut[27][8];
              muxOutConnector[44] = fifoOut[28][8];
              muxOutConnector[45] = fifoOut[29][8];
              muxOutConnector[46] = fifoOut[30][8];
              muxOutConnector[47] = fifoOut[31][8];
              muxOutConnector[48] = fifoOut[32][8];
              muxOutConnector[49] = fifoOut[33][8];
              muxOutConnector[50] = fifoOut[34][8];
              muxOutConnector[51] = fifoOut[35][8];
         end
         17: begin
              muxOutConnector[0] = fifoOut[8][6];
              muxOutConnector[1] = fifoOut[9][6];
              muxOutConnector[2] = fifoOut[10][6];
              muxOutConnector[3] = fifoOut[11][6];
              muxOutConnector[4] = fifoOut[12][6];
              muxOutConnector[5] = fifoOut[13][6];
              muxOutConnector[6] = fifoOut[14][6];
              muxOutConnector[7] = fifoOut[15][6];
              muxOutConnector[8] = fifoOut[16][6];
              muxOutConnector[9] = fifoOut[17][6];
              muxOutConnector[10] = fifoOut[18][6];
              muxOutConnector[11] = fifoOut[19][6];
              muxOutConnector[12] = fifoOut[20][6];
              muxOutConnector[13] = fifoOut[21][6];
              muxOutConnector[14] = fifoOut[22][6];
              muxOutConnector[15] = fifoOut[23][6];
              muxOutConnector[16] = fifoOut[24][6];
              muxOutConnector[17] = fifoOut[25][6];
              muxOutConnector[18] = fifoOut[0][5];
              muxOutConnector[19] = fifoOut[1][5];
              muxOutConnector[20] = fifoOut[2][5];
              muxOutConnector[21] = fifoOut[3][5];
              muxOutConnector[22] = fifoOut[4][5];
              muxOutConnector[23] = fifoOut[5][5];
              muxOutConnector[24] = fifoOut[6][5];
              muxOutConnector[25] = fifoOut[7][5];
              muxOutConnector[26] = fifoOut[36][9];
              muxOutConnector[27] = fifoOut[37][9];
              muxOutConnector[28] = fifoOut[38][9];
              muxOutConnector[29] = fifoOut[39][9];
              muxOutConnector[30] = fifoOut[40][9];
              muxOutConnector[31] = fifoOut[41][9];
              muxOutConnector[32] = fifoOut[42][9];
              muxOutConnector[33] = fifoOut[43][9];
              muxOutConnector[34] = fifoOut[44][9];
              muxOutConnector[35] = fifoOut[45][9];
              muxOutConnector[36] = fifoOut[46][9];
              muxOutConnector[37] = fifoOut[47][9];
              muxOutConnector[38] = fifoOut[48][9];
              muxOutConnector[39] = fifoOut[49][9];
              muxOutConnector[40] = fifoOut[50][9];
              muxOutConnector[41] = fifoOut[51][9];
              muxOutConnector[42] = fifoOut[26][8];
              muxOutConnector[43] = fifoOut[27][8];
              muxOutConnector[44] = fifoOut[28][8];
              muxOutConnector[45] = fifoOut[29][8];
              muxOutConnector[46] = fifoOut[30][8];
              muxOutConnector[47] = fifoOut[31][8];
              muxOutConnector[48] = fifoOut[32][8];
              muxOutConnector[49] = fifoOut[33][8];
              muxOutConnector[50] = fifoOut[34][8];
              muxOutConnector[51] = fifoOut[35][8];
         end
         18: begin
              muxOutConnector[0] = fifoOut[8][6];
              muxOutConnector[1] = fifoOut[9][6];
              muxOutConnector[2] = fifoOut[10][6];
              muxOutConnector[3] = fifoOut[11][6];
              muxOutConnector[4] = fifoOut[12][6];
              muxOutConnector[5] = fifoOut[13][6];
              muxOutConnector[6] = fifoOut[14][6];
              muxOutConnector[7] = fifoOut[15][6];
              muxOutConnector[8] = fifoOut[16][6];
              muxOutConnector[9] = fifoOut[17][6];
              muxOutConnector[10] = fifoOut[18][6];
              muxOutConnector[11] = fifoOut[19][6];
              muxOutConnector[12] = fifoOut[20][6];
              muxOutConnector[13] = fifoOut[21][6];
              muxOutConnector[14] = fifoOut[22][6];
              muxOutConnector[15] = fifoOut[23][6];
              muxOutConnector[16] = fifoOut[24][6];
              muxOutConnector[17] = fifoOut[25][6];
              muxOutConnector[18] = fifoOut[0][5];
              muxOutConnector[19] = fifoOut[1][5];
              muxOutConnector[20] = fifoOut[2][5];
              muxOutConnector[21] = fifoOut[3][5];
              muxOutConnector[22] = fifoOut[4][5];
              muxOutConnector[23] = fifoOut[5][5];
              muxOutConnector[24] = fifoOut[6][5];
              muxOutConnector[25] = fifoOut[7][5];
              muxOutConnector[26] = fifoOut[36][9];
              muxOutConnector[27] = fifoOut[37][9];
              muxOutConnector[28] = fifoOut[38][9];
              muxOutConnector[29] = fifoOut[39][9];
              muxOutConnector[30] = fifoOut[40][9];
              muxOutConnector[31] = fifoOut[41][9];
              muxOutConnector[32] = fifoOut[42][9];
              muxOutConnector[33] = fifoOut[43][9];
              muxOutConnector[34] = fifoOut[44][9];
              muxOutConnector[35] = fifoOut[45][9];
              muxOutConnector[36] = fifoOut[46][9];
              muxOutConnector[37] = fifoOut[47][9];
              muxOutConnector[38] = fifoOut[48][9];
              muxOutConnector[39] = fifoOut[49][9];
              muxOutConnector[40] = fifoOut[50][9];
              muxOutConnector[41] = fifoOut[51][9];
              muxOutConnector[42] = fifoOut[26][8];
              muxOutConnector[43] = fifoOut[27][8];
              muxOutConnector[44] = fifoOut[28][8];
              muxOutConnector[45] = fifoOut[29][8];
              muxOutConnector[46] = fifoOut[30][8];
              muxOutConnector[47] = fifoOut[31][8];
              muxOutConnector[48] = fifoOut[32][8];
              muxOutConnector[49] = fifoOut[33][8];
              muxOutConnector[50] = fifoOut[34][8];
              muxOutConnector[51] = fifoOut[35][8];
         end
         19: begin
              muxOutConnector[0] = fifoOut[8][6];
              muxOutConnector[1] = fifoOut[9][6];
              muxOutConnector[2] = fifoOut[10][6];
              muxOutConnector[3] = fifoOut[11][6];
              muxOutConnector[4] = fifoOut[12][6];
              muxOutConnector[5] = fifoOut[13][6];
              muxOutConnector[6] = fifoOut[14][6];
              muxOutConnector[7] = fifoOut[15][6];
              muxOutConnector[8] = fifoOut[16][6];
              muxOutConnector[9] = fifoOut[17][6];
              muxOutConnector[10] = fifoOut[18][6];
              muxOutConnector[11] = fifoOut[19][6];
              muxOutConnector[12] = fifoOut[20][6];
              muxOutConnector[13] = fifoOut[21][6];
              muxOutConnector[14] = fifoOut[22][6];
              muxOutConnector[15] = fifoOut[23][6];
              muxOutConnector[16] = fifoOut[24][6];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[36][9];
              muxOutConnector[27] = fifoOut[37][9];
              muxOutConnector[28] = fifoOut[38][9];
              muxOutConnector[29] = fifoOut[39][9];
              muxOutConnector[30] = fifoOut[40][9];
              muxOutConnector[31] = fifoOut[41][9];
              muxOutConnector[32] = fifoOut[42][9];
              muxOutConnector[33] = fifoOut[43][9];
              muxOutConnector[34] = fifoOut[44][9];
              muxOutConnector[35] = fifoOut[45][9];
              muxOutConnector[36] = fifoOut[46][9];
              muxOutConnector[37] = fifoOut[47][9];
              muxOutConnector[38] = fifoOut[48][9];
              muxOutConnector[39] = fifoOut[49][9];
              muxOutConnector[40] = fifoOut[50][9];
              muxOutConnector[41] = fifoOut[51][9];
              muxOutConnector[42] = fifoOut[26][8];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
         end
         default: begin
               for(i=0;i<muxOutSymbols;i=i+1)begin
                muxOutConnector[i] = 0;
              end
         end
//hgjhgbuiguigbigbgbgbui
         endcase
         end
         endcase
         end
endmodule