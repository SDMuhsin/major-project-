`timescale 1ns / 1ps
module LMem1To0_511_circ4_combined_ns_yu_pipelined_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        rxIn,
        load_input_en,
        iteration_0_indicator,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter r_lower = 32;
parameter c = 17;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input [ADDRESSWIDTH-1:0]unloadAddress;
input load_input_en;
input iteration_0_indicator;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input [ r_lower * w - 1 : 0 ] rxIn; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
reg [ w - 1 : 0 ]column_1[ r - 1 : 0 ];
reg chip_en;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
wire [w-1:0]rxInConnector[r_lower-1:0]; // Change #
reg [ muxOutSymbols * w - 1 : 0]muxOut_firstiter_reg0, muxOut_process_reg0;
wire [ muxOutSymbols * w - 1 : 0]muxOut_firstiter, muxOut_process;
reg [w-1:0]muxOutConnector_firstiter[ muxOutSymbols  - 1 : 0];
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

 assign muxOut = iteration_0_indicator ? muxOut_firstiter_reg0 : muxOut_process_reg0;
always@(posedge clk)begin
    if (!rst) begin
      muxOut_firstiter_reg0 <= 0;
      muxOut_process_reg0 <= 0;
    end
    else begin
      muxOut_firstiter_reg0 <= muxOut_firstiter;
      muxOut_process_reg0 <= muxOut_process;
    end
end

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut_firstiter[ (k+1)*w-1:k*w] = muxOutConnector_firstiter[k];
        assign muxOut_process[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

generate
    for (k=0;k<r_lower;k=k+1)begin:assign_rx
        assign rxInConnector[k] = rxIn[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (!rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(chip_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            fifoOut[i][0] <= column_1[i];
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

    always@(*) begin
      if(load_input_en)begin
        chip_en=load_input_en;
      end
      else if(wr_en)begin
        chip_en=wr_en;
      end
      else begin // if wr_en or load_en=0, dont shift or load inputs
        chip_en=0;
      end
      for(i = r-1; i > -1; i=i-1) begin
        if(load_input_en)begin
          if(i < r_lower)begin
             column_1[i] = rxInConnector[i];
          end
          else begin
             column_1[i] = maxVal;
          end
        end
        else begin//wr_en=1 or 0 or load_en=0 case: connect input but loading does not happen since chipen=0
          column_1[i] <= ly0InConnector[i];
        end
      end
    end//always
assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
       0: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = fifoOut[10][8][w-1];
              unloadMuxOut[11] = fifoOut[11][8][w-1];
              unloadMuxOut[12] = fifoOut[12][8][w-1];
              unloadMuxOut[13] = fifoOut[13][8][w-1];
              unloadMuxOut[14] = fifoOut[14][8][w-1];
              unloadMuxOut[15] = fifoOut[15][8][w-1];
              unloadMuxOut[16] = fifoOut[16][8][w-1];
              unloadMuxOut[17] = fifoOut[17][8][w-1];
              unloadMuxOut[18] = fifoOut[18][8][w-1];
              unloadMuxOut[19] = fifoOut[19][8][w-1];
              unloadMuxOut[20] = fifoOut[20][8][w-1];
              unloadMuxOut[21] = fifoOut[21][8][w-1];
              unloadMuxOut[22] = fifoOut[22][8][w-1];
              unloadMuxOut[23] = fifoOut[23][8][w-1];
              unloadMuxOut[24] = fifoOut[24][8][w-1];
              unloadMuxOut[25] = fifoOut[25][8][w-1];
              unloadMuxOut[26] = fifoOut[0][7][w-1];
              unloadMuxOut[27] = fifoOut[1][7][w-1];
              unloadMuxOut[28] = fifoOut[2][7][w-1];
              unloadMuxOut[29] = fifoOut[3][7][w-1];
              unloadMuxOut[30] = fifoOut[4][7][w-1];
              unloadMuxOut[31] = fifoOut[5][7][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[6][7][w-1];
              unloadMuxOut[1] = fifoOut[7][7][w-1];
              unloadMuxOut[2] = fifoOut[8][7][w-1];
              unloadMuxOut[3] = fifoOut[9][7][w-1];
              unloadMuxOut[4] = fifoOut[10][7][w-1];
              unloadMuxOut[5] = fifoOut[11][7][w-1];
              unloadMuxOut[6] = fifoOut[12][7][w-1];
              unloadMuxOut[7] = fifoOut[13][7][w-1];
              unloadMuxOut[8] = fifoOut[14][7][w-1];
              unloadMuxOut[9] = fifoOut[15][7][w-1];
              unloadMuxOut[10] = fifoOut[16][7][w-1];
              unloadMuxOut[11] = fifoOut[17][7][w-1];
              unloadMuxOut[12] = fifoOut[18][7][w-1];
              unloadMuxOut[13] = fifoOut[19][7][w-1];
              unloadMuxOut[14] = fifoOut[20][7][w-1];
              unloadMuxOut[15] = fifoOut[21][7][w-1];
              unloadMuxOut[16] = fifoOut[22][7][w-1];
              unloadMuxOut[17] = fifoOut[23][7][w-1];
              unloadMuxOut[18] = fifoOut[24][7][w-1];
              unloadMuxOut[19] = fifoOut[25][7][w-1];
              unloadMuxOut[20] = fifoOut[0][6][w-1];
              unloadMuxOut[21] = fifoOut[1][6][w-1];
              unloadMuxOut[22] = fifoOut[2][6][w-1];
              unloadMuxOut[23] = fifoOut[3][6][w-1];
              unloadMuxOut[24] = fifoOut[4][6][w-1];
              unloadMuxOut[25] = fifoOut[5][6][w-1];
              unloadMuxOut[26] = fifoOut[6][6][w-1];
              unloadMuxOut[27] = fifoOut[7][6][w-1];
              unloadMuxOut[28] = fifoOut[8][6][w-1];
              unloadMuxOut[29] = fifoOut[9][6][w-1];
              unloadMuxOut[30] = fifoOut[10][6][w-1];
              unloadMuxOut[31] = fifoOut[11][6][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[12][6][w-1];
              unloadMuxOut[1] = fifoOut[13][6][w-1];
              unloadMuxOut[2] = fifoOut[14][6][w-1];
              unloadMuxOut[3] = fifoOut[15][6][w-1];
              unloadMuxOut[4] = fifoOut[16][6][w-1];
              unloadMuxOut[5] = fifoOut[17][6][w-1];
              unloadMuxOut[6] = fifoOut[18][6][w-1];
              unloadMuxOut[7] = fifoOut[19][6][w-1];
              unloadMuxOut[8] = fifoOut[20][6][w-1];
              unloadMuxOut[9] = fifoOut[21][6][w-1];
              unloadMuxOut[10] = fifoOut[22][6][w-1];
              unloadMuxOut[11] = fifoOut[23][6][w-1];
              unloadMuxOut[12] = fifoOut[24][6][w-1];
              unloadMuxOut[13] = fifoOut[25][6][w-1];
              unloadMuxOut[14] = fifoOut[0][5][w-1];
              unloadMuxOut[15] = fifoOut[1][5][w-1];
              unloadMuxOut[16] = fifoOut[2][5][w-1];
              unloadMuxOut[17] = fifoOut[3][5][w-1];
              unloadMuxOut[18] = fifoOut[4][5][w-1];
              unloadMuxOut[19] = fifoOut[5][5][w-1];
              unloadMuxOut[20] = fifoOut[6][5][w-1];
              unloadMuxOut[21] = fifoOut[7][5][w-1];
              unloadMuxOut[22] = fifoOut[8][5][w-1];
              unloadMuxOut[23] = fifoOut[9][5][w-1];
              unloadMuxOut[24] = fifoOut[10][5][w-1];
              unloadMuxOut[25] = fifoOut[11][5][w-1];
              unloadMuxOut[26] = fifoOut[12][5][w-1];
              unloadMuxOut[27] = fifoOut[13][5][w-1];
              unloadMuxOut[28] = fifoOut[14][5][w-1];
              unloadMuxOut[29] = fifoOut[15][5][w-1];
              unloadMuxOut[30] = fifoOut[16][5][w-1];
              unloadMuxOut[31] = fifoOut[17][5][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[18][5][w-1];
              unloadMuxOut[1] = fifoOut[19][5][w-1];
              unloadMuxOut[2] = fifoOut[20][5][w-1];
              unloadMuxOut[3] = fifoOut[21][5][w-1];
              unloadMuxOut[4] = fifoOut[22][5][w-1];
              unloadMuxOut[5] = fifoOut[23][5][w-1];
              unloadMuxOut[6] = fifoOut[24][5][w-1];
              unloadMuxOut[7] = fifoOut[25][5][w-1];
              unloadMuxOut[8] = fifoOut[0][4][w-1];
              unloadMuxOut[9] = fifoOut[1][4][w-1];
              unloadMuxOut[10] = fifoOut[2][4][w-1];
              unloadMuxOut[11] = fifoOut[3][4][w-1];
              unloadMuxOut[12] = fifoOut[4][4][w-1];
              unloadMuxOut[13] = fifoOut[5][4][w-1];
              unloadMuxOut[14] = fifoOut[6][4][w-1];
              unloadMuxOut[15] = fifoOut[7][4][w-1];
              unloadMuxOut[16] = fifoOut[8][4][w-1];
              unloadMuxOut[17] = fifoOut[9][4][w-1];
              unloadMuxOut[18] = fifoOut[10][4][w-1];
              unloadMuxOut[19] = fifoOut[11][4][w-1];
              unloadMuxOut[20] = fifoOut[12][4][w-1];
              unloadMuxOut[21] = fifoOut[13][4][w-1];
              unloadMuxOut[22] = fifoOut[14][4][w-1];
              unloadMuxOut[23] = fifoOut[15][4][w-1];
              unloadMuxOut[24] = fifoOut[16][4][w-1];
              unloadMuxOut[25] = fifoOut[17][4][w-1];
              unloadMuxOut[26] = fifoOut[18][4][w-1];
              unloadMuxOut[27] = fifoOut[19][4][w-1];
              unloadMuxOut[28] = fifoOut[20][4][w-1];
              unloadMuxOut[29] = fifoOut[21][4][w-1];
              unloadMuxOut[30] = fifoOut[22][4][w-1];
              unloadMuxOut[31] = fifoOut[23][4][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[24][4][w-1];
              unloadMuxOut[1] = fifoOut[25][4][w-1];
              unloadMuxOut[2] = fifoOut[0][3][w-1];
              unloadMuxOut[3] = fifoOut[1][3][w-1];
              unloadMuxOut[4] = fifoOut[2][3][w-1];
              unloadMuxOut[5] = fifoOut[3][3][w-1];
              unloadMuxOut[6] = fifoOut[4][3][w-1];
              unloadMuxOut[7] = fifoOut[5][3][w-1];
              unloadMuxOut[8] = fifoOut[6][3][w-1];
              unloadMuxOut[9] = fifoOut[7][3][w-1];
              unloadMuxOut[10] = fifoOut[8][3][w-1];
              unloadMuxOut[11] = fifoOut[9][3][w-1];
              unloadMuxOut[12] = fifoOut[10][3][w-1];
              unloadMuxOut[13] = fifoOut[11][3][w-1];
              unloadMuxOut[14] = fifoOut[12][3][w-1];
              unloadMuxOut[15] = fifoOut[13][3][w-1];
              unloadMuxOut[16] = fifoOut[14][3][w-1];
              unloadMuxOut[17] = fifoOut[15][3][w-1];
              unloadMuxOut[18] = fifoOut[16][3][w-1];
              unloadMuxOut[19] = fifoOut[17][3][w-1];
              unloadMuxOut[20] = fifoOut[18][3][w-1];
              unloadMuxOut[21] = fifoOut[19][3][w-1];
              unloadMuxOut[22] = fifoOut[20][3][w-1];
              unloadMuxOut[23] = fifoOut[21][3][w-1];
              unloadMuxOut[24] = fifoOut[22][3][w-1];
              unloadMuxOut[25] = fifoOut[23][3][w-1];
              unloadMuxOut[26] = fifoOut[24][3][w-1];
              unloadMuxOut[27] = fifoOut[25][3][w-1];
              unloadMuxOut[28] = fifoOut[0][2][w-1];
              unloadMuxOut[29] = fifoOut[1][2][w-1];
              unloadMuxOut[30] = fifoOut[2][2][w-1];
              unloadMuxOut[31] = fifoOut[3][2][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[4][2][w-1];
              unloadMuxOut[1] = fifoOut[5][2][w-1];
              unloadMuxOut[2] = fifoOut[6][2][w-1];
              unloadMuxOut[3] = fifoOut[7][2][w-1];
              unloadMuxOut[4] = fifoOut[8][2][w-1];
              unloadMuxOut[5] = fifoOut[9][2][w-1];
              unloadMuxOut[6] = fifoOut[10][2][w-1];
              unloadMuxOut[7] = fifoOut[11][2][w-1];
              unloadMuxOut[8] = fifoOut[12][2][w-1];
              unloadMuxOut[9] = fifoOut[13][2][w-1];
              unloadMuxOut[10] = fifoOut[14][2][w-1];
              unloadMuxOut[11] = fifoOut[15][2][w-1];
              unloadMuxOut[12] = fifoOut[16][2][w-1];
              unloadMuxOut[13] = fifoOut[17][2][w-1];
              unloadMuxOut[14] = fifoOut[18][2][w-1];
              unloadMuxOut[15] = fifoOut[19][2][w-1];
              unloadMuxOut[16] = fifoOut[20][2][w-1];
              unloadMuxOut[17] = fifoOut[21][2][w-1];
              unloadMuxOut[18] = fifoOut[22][2][w-1];
              unloadMuxOut[19] = fifoOut[23][2][w-1];
              unloadMuxOut[20] = fifoOut[24][2][w-1];
              unloadMuxOut[21] = fifoOut[25][2][w-1];
              unloadMuxOut[22] = fifoOut[0][1][w-1];
              unloadMuxOut[23] = fifoOut[1][1][w-1];
              unloadMuxOut[24] = fifoOut[2][1][w-1];
              unloadMuxOut[25] = fifoOut[3][1][w-1];
              unloadMuxOut[26] = fifoOut[4][1][w-1];
              unloadMuxOut[27] = fifoOut[5][1][w-1];
              unloadMuxOut[28] = fifoOut[6][1][w-1];
              unloadMuxOut[29] = fifoOut[7][1][w-1];
              unloadMuxOut[30] = fifoOut[8][1][w-1];
              unloadMuxOut[31] = fifoOut[9][1][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[10][1][w-1];
              unloadMuxOut[1] = fifoOut[11][1][w-1];
              unloadMuxOut[2] = fifoOut[12][1][w-1];
              unloadMuxOut[3] = fifoOut[13][1][w-1];
              unloadMuxOut[4] = fifoOut[14][1][w-1];
              unloadMuxOut[5] = fifoOut[15][1][w-1];
              unloadMuxOut[6] = fifoOut[16][1][w-1];
              unloadMuxOut[7] = fifoOut[17][1][w-1];
              unloadMuxOut[8] = fifoOut[18][1][w-1];
              unloadMuxOut[9] = fifoOut[19][1][w-1];
              unloadMuxOut[10] = fifoOut[20][1][w-1];
              unloadMuxOut[11] = fifoOut[21][1][w-1];
              unloadMuxOut[12] = fifoOut[22][1][w-1];
              unloadMuxOut[13] = fifoOut[23][1][w-1];
              unloadMuxOut[14] = fifoOut[24][1][w-1];
              unloadMuxOut[15] = fifoOut[25][1][w-1];
              unloadMuxOut[16] = fifoOut[0][0][w-1];
              unloadMuxOut[17] = fifoOut[1][0][w-1];
              unloadMuxOut[18] = fifoOut[2][0][w-1];
              unloadMuxOut[19] = fifoOut[3][0][w-1];
              unloadMuxOut[20] = fifoOut[4][0][w-1];
              unloadMuxOut[21] = fifoOut[5][0][w-1];
              unloadMuxOut[22] = fifoOut[6][0][w-1];
              unloadMuxOut[23] = fifoOut[7][0][w-1];
              unloadMuxOut[24] = fifoOut[8][0][w-1];
              unloadMuxOut[25] = fifoOut[9][0][w-1];
              unloadMuxOut[26] = fifoOut[10][0][w-1];
              unloadMuxOut[27] = fifoOut[11][0][w-1];
              unloadMuxOut[28] = fifoOut[12][0][w-1];
              unloadMuxOut[29] = fifoOut[13][0][w-1];
              unloadMuxOut[30] = fifoOut[14][0][w-1];
              unloadMuxOut[31] = fifoOut[15][0][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[16][0][w-1];
              unloadMuxOut[1] = fifoOut[46][8][w-1];
              unloadMuxOut[2] = fifoOut[47][8][w-1];
              unloadMuxOut[3] = fifoOut[48][8][w-1];
              unloadMuxOut[4] = fifoOut[49][8][w-1];
              unloadMuxOut[5] = fifoOut[50][8][w-1];
              unloadMuxOut[6] = fifoOut[51][8][w-1];
              unloadMuxOut[7] = fifoOut[26][7][w-1];
              unloadMuxOut[8] = fifoOut[27][7][w-1];
              unloadMuxOut[9] = fifoOut[28][7][w-1];
              unloadMuxOut[10] = fifoOut[29][7][w-1];
              unloadMuxOut[11] = fifoOut[30][7][w-1];
              unloadMuxOut[12] = fifoOut[31][7][w-1];
              unloadMuxOut[13] = fifoOut[32][7][w-1];
              unloadMuxOut[14] = fifoOut[33][7][w-1];
              unloadMuxOut[15] = fifoOut[34][7][w-1];
              unloadMuxOut[16] = fifoOut[35][7][w-1];
              unloadMuxOut[17] = fifoOut[36][7][w-1];
              unloadMuxOut[18] = fifoOut[37][7][w-1];
              unloadMuxOut[19] = fifoOut[38][7][w-1];
              unloadMuxOut[20] = fifoOut[39][7][w-1];
              unloadMuxOut[21] = fifoOut[40][7][w-1];
              unloadMuxOut[22] = fifoOut[41][7][w-1];
              unloadMuxOut[23] = fifoOut[42][7][w-1];
              unloadMuxOut[24] = fifoOut[43][7][w-1];
              unloadMuxOut[25] = fifoOut[44][7][w-1];
              unloadMuxOut[26] = fifoOut[45][7][w-1];
              unloadMuxOut[27] = fifoOut[46][7][w-1];
              unloadMuxOut[28] = fifoOut[47][7][w-1];
              unloadMuxOut[29] = fifoOut[48][7][w-1];
              unloadMuxOut[30] = fifoOut[49][7][w-1];
              unloadMuxOut[31] = fifoOut[50][7][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[51][7][w-1];
              unloadMuxOut[1] = fifoOut[26][6][w-1];
              unloadMuxOut[2] = fifoOut[27][6][w-1];
              unloadMuxOut[3] = fifoOut[28][6][w-1];
              unloadMuxOut[4] = fifoOut[29][6][w-1];
              unloadMuxOut[5] = fifoOut[30][6][w-1];
              unloadMuxOut[6] = fifoOut[31][6][w-1];
              unloadMuxOut[7] = fifoOut[32][6][w-1];
              unloadMuxOut[8] = fifoOut[33][6][w-1];
              unloadMuxOut[9] = fifoOut[34][6][w-1];
              unloadMuxOut[10] = fifoOut[35][6][w-1];
              unloadMuxOut[11] = fifoOut[36][6][w-1];
              unloadMuxOut[12] = fifoOut[37][6][w-1];
              unloadMuxOut[13] = fifoOut[38][6][w-1];
              unloadMuxOut[14] = fifoOut[39][6][w-1];
              unloadMuxOut[15] = fifoOut[40][6][w-1];
              unloadMuxOut[16] = fifoOut[41][6][w-1];
              unloadMuxOut[17] = fifoOut[42][6][w-1];
              unloadMuxOut[18] = fifoOut[43][6][w-1];
              unloadMuxOut[19] = fifoOut[44][6][w-1];
              unloadMuxOut[20] = fifoOut[45][6][w-1];
              unloadMuxOut[21] = fifoOut[46][6][w-1];
              unloadMuxOut[22] = fifoOut[47][6][w-1];
              unloadMuxOut[23] = fifoOut[48][6][w-1];
              unloadMuxOut[24] = fifoOut[49][6][w-1];
              unloadMuxOut[25] = fifoOut[50][6][w-1];
              unloadMuxOut[26] = fifoOut[51][6][w-1];
              unloadMuxOut[27] = fifoOut[26][5][w-1];
              unloadMuxOut[28] = fifoOut[27][5][w-1];
              unloadMuxOut[29] = fifoOut[28][5][w-1];
              unloadMuxOut[30] = fifoOut[29][5][w-1];
              unloadMuxOut[31] = fifoOut[30][5][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[31][5][w-1];
              unloadMuxOut[1] = fifoOut[32][5][w-1];
              unloadMuxOut[2] = fifoOut[33][5][w-1];
              unloadMuxOut[3] = fifoOut[34][5][w-1];
              unloadMuxOut[4] = fifoOut[35][5][w-1];
              unloadMuxOut[5] = fifoOut[36][5][w-1];
              unloadMuxOut[6] = fifoOut[37][5][w-1];
              unloadMuxOut[7] = fifoOut[38][5][w-1];
              unloadMuxOut[8] = fifoOut[39][5][w-1];
              unloadMuxOut[9] = fifoOut[40][5][w-1];
              unloadMuxOut[10] = fifoOut[41][5][w-1];
              unloadMuxOut[11] = fifoOut[42][5][w-1];
              unloadMuxOut[12] = fifoOut[43][5][w-1];
              unloadMuxOut[13] = fifoOut[44][5][w-1];
              unloadMuxOut[14] = fifoOut[45][5][w-1];
              unloadMuxOut[15] = fifoOut[46][5][w-1];
              unloadMuxOut[16] = fifoOut[47][5][w-1];
              unloadMuxOut[17] = fifoOut[48][5][w-1];
              unloadMuxOut[18] = fifoOut[49][5][w-1];
              unloadMuxOut[19] = fifoOut[50][5][w-1];
              unloadMuxOut[20] = fifoOut[51][5][w-1];
              unloadMuxOut[21] = fifoOut[26][4][w-1];
              unloadMuxOut[22] = fifoOut[27][4][w-1];
              unloadMuxOut[23] = fifoOut[28][4][w-1];
              unloadMuxOut[24] = fifoOut[29][4][w-1];
              unloadMuxOut[25] = fifoOut[30][4][w-1];
              unloadMuxOut[26] = fifoOut[31][4][w-1];
              unloadMuxOut[27] = fifoOut[32][4][w-1];
              unloadMuxOut[28] = fifoOut[33][4][w-1];
              unloadMuxOut[29] = fifoOut[34][4][w-1];
              unloadMuxOut[30] = fifoOut[35][4][w-1];
              unloadMuxOut[31] = fifoOut[36][4][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[37][4][w-1];
              unloadMuxOut[1] = fifoOut[38][4][w-1];
              unloadMuxOut[2] = fifoOut[39][4][w-1];
              unloadMuxOut[3] = fifoOut[40][4][w-1];
              unloadMuxOut[4] = fifoOut[41][4][w-1];
              unloadMuxOut[5] = fifoOut[42][4][w-1];
              unloadMuxOut[6] = fifoOut[43][4][w-1];
              unloadMuxOut[7] = fifoOut[44][4][w-1];
              unloadMuxOut[8] = fifoOut[45][4][w-1];
              unloadMuxOut[9] = fifoOut[46][4][w-1];
              unloadMuxOut[10] = fifoOut[47][4][w-1];
              unloadMuxOut[11] = fifoOut[48][4][w-1];
              unloadMuxOut[12] = fifoOut[49][4][w-1];
              unloadMuxOut[13] = fifoOut[50][4][w-1];
              unloadMuxOut[14] = fifoOut[51][4][w-1];
              unloadMuxOut[15] = fifoOut[26][3][w-1];
              unloadMuxOut[16] = fifoOut[27][3][w-1];
              unloadMuxOut[17] = fifoOut[28][3][w-1];
              unloadMuxOut[18] = fifoOut[29][3][w-1];
              unloadMuxOut[19] = fifoOut[30][3][w-1];
              unloadMuxOut[20] = fifoOut[31][3][w-1];
              unloadMuxOut[21] = fifoOut[32][3][w-1];
              unloadMuxOut[22] = fifoOut[33][3][w-1];
              unloadMuxOut[23] = fifoOut[34][3][w-1];
              unloadMuxOut[24] = fifoOut[35][3][w-1];
              unloadMuxOut[25] = fifoOut[36][3][w-1];
              unloadMuxOut[26] = fifoOut[37][3][w-1];
              unloadMuxOut[27] = fifoOut[38][3][w-1];
              unloadMuxOut[28] = fifoOut[39][3][w-1];
              unloadMuxOut[29] = fifoOut[40][3][w-1];
              unloadMuxOut[30] = fifoOut[41][3][w-1];
              unloadMuxOut[31] = fifoOut[42][3][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[43][3][w-1];
              unloadMuxOut[1] = fifoOut[44][3][w-1];
              unloadMuxOut[2] = fifoOut[45][3][w-1];
              unloadMuxOut[3] = fifoOut[46][3][w-1];
              unloadMuxOut[4] = fifoOut[47][3][w-1];
              unloadMuxOut[5] = fifoOut[48][3][w-1];
              unloadMuxOut[6] = fifoOut[49][3][w-1];
              unloadMuxOut[7] = fifoOut[50][3][w-1];
              unloadMuxOut[8] = fifoOut[51][3][w-1];
              unloadMuxOut[9] = fifoOut[26][2][w-1];
              unloadMuxOut[10] = fifoOut[27][2][w-1];
              unloadMuxOut[11] = fifoOut[28][2][w-1];
              unloadMuxOut[12] = fifoOut[29][2][w-1];
              unloadMuxOut[13] = fifoOut[30][2][w-1];
              unloadMuxOut[14] = fifoOut[31][2][w-1];
              unloadMuxOut[15] = fifoOut[32][2][w-1];
              unloadMuxOut[16] = fifoOut[33][2][w-1];
              unloadMuxOut[17] = fifoOut[34][2][w-1];
              unloadMuxOut[18] = fifoOut[35][2][w-1];
              unloadMuxOut[19] = fifoOut[36][2][w-1];
              unloadMuxOut[20] = fifoOut[37][2][w-1];
              unloadMuxOut[21] = fifoOut[38][2][w-1];
              unloadMuxOut[22] = fifoOut[39][2][w-1];
              unloadMuxOut[23] = fifoOut[40][2][w-1];
              unloadMuxOut[24] = fifoOut[41][2][w-1];
              unloadMuxOut[25] = fifoOut[42][2][w-1];
              unloadMuxOut[26] = fifoOut[43][2][w-1];
              unloadMuxOut[27] = fifoOut[44][2][w-1];
              unloadMuxOut[28] = fifoOut[45][2][w-1];
              unloadMuxOut[29] = fifoOut[46][2][w-1];
              unloadMuxOut[30] = fifoOut[47][2][w-1];
              unloadMuxOut[31] = fifoOut[48][2][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[49][2][w-1];
              unloadMuxOut[1] = fifoOut[50][2][w-1];
              unloadMuxOut[2] = fifoOut[51][2][w-1];
              unloadMuxOut[3] = fifoOut[26][1][w-1];
              unloadMuxOut[4] = fifoOut[27][1][w-1];
              unloadMuxOut[5] = fifoOut[28][1][w-1];
              unloadMuxOut[6] = fifoOut[29][1][w-1];
              unloadMuxOut[7] = fifoOut[30][1][w-1];
              unloadMuxOut[8] = fifoOut[31][1][w-1];
              unloadMuxOut[9] = fifoOut[32][1][w-1];
              unloadMuxOut[10] = fifoOut[33][1][w-1];
              unloadMuxOut[11] = fifoOut[34][1][w-1];
              unloadMuxOut[12] = fifoOut[35][1][w-1];
              unloadMuxOut[13] = fifoOut[36][1][w-1];
              unloadMuxOut[14] = fifoOut[37][1][w-1];
              unloadMuxOut[15] = fifoOut[38][1][w-1];
              unloadMuxOut[16] = fifoOut[39][1][w-1];
              unloadMuxOut[17] = fifoOut[40][1][w-1];
              unloadMuxOut[18] = fifoOut[41][1][w-1];
              unloadMuxOut[19] = fifoOut[42][1][w-1];
              unloadMuxOut[20] = fifoOut[43][1][w-1];
              unloadMuxOut[21] = fifoOut[44][1][w-1];
              unloadMuxOut[22] = fifoOut[45][1][w-1];
              unloadMuxOut[23] = fifoOut[46][1][w-1];
              unloadMuxOut[24] = fifoOut[47][1][w-1];
              unloadMuxOut[25] = fifoOut[48][1][w-1];
              unloadMuxOut[26] = fifoOut[49][1][w-1];
              unloadMuxOut[27] = fifoOut[50][1][w-1];
              unloadMuxOut[28] = fifoOut[51][1][w-1];
              unloadMuxOut[29] = fifoOut[26][0][w-1];
              unloadMuxOut[30] = fifoOut[27][0][w-1];
              unloadMuxOut[31] = fifoOut[28][0][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[29][0][w-1];
              unloadMuxOut[1] = fifoOut[30][0][w-1];
              unloadMuxOut[2] = fifoOut[31][0][w-1];
              unloadMuxOut[3] = fifoOut[32][0][w-1];
              unloadMuxOut[4] = fifoOut[33][0][w-1];
              unloadMuxOut[5] = fifoOut[34][0][w-1];
              unloadMuxOut[6] = fifoOut[35][0][w-1];
              unloadMuxOut[7] = fifoOut[36][0][w-1];
              unloadMuxOut[8] = fifoOut[37][0][w-1];
              unloadMuxOut[9] = fifoOut[38][0][w-1];
              unloadMuxOut[10] = fifoOut[39][0][w-1];
              unloadMuxOut[11] = fifoOut[40][0][w-1];
              unloadMuxOut[12] = fifoOut[41][0][w-1];
              unloadMuxOut[13] = fifoOut[42][0][w-1];
              unloadMuxOut[14] = fifoOut[23][12][w-1];
              unloadMuxOut[15] = fifoOut[24][12][w-1];
              unloadMuxOut[16] = fifoOut[25][12][w-1];
              unloadMuxOut[17] = fifoOut[0][11][w-1];
              unloadMuxOut[18] = fifoOut[1][11][w-1];
              unloadMuxOut[19] = fifoOut[2][11][w-1];
              unloadMuxOut[20] = fifoOut[3][11][w-1];
              unloadMuxOut[21] = fifoOut[4][11][w-1];
              unloadMuxOut[22] = fifoOut[5][11][w-1];
              unloadMuxOut[23] = fifoOut[6][11][w-1];
              unloadMuxOut[24] = fifoOut[7][11][w-1];
              unloadMuxOut[25] = fifoOut[8][11][w-1];
              unloadMuxOut[26] = fifoOut[9][11][w-1];
              unloadMuxOut[27] = fifoOut[10][11][w-1];
              unloadMuxOut[28] = fifoOut[11][11][w-1];
              unloadMuxOut[29] = fifoOut[12][11][w-1];
              unloadMuxOut[30] = fifoOut[13][11][w-1];
              unloadMuxOut[31] = fifoOut[14][11][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[15][11][w-1];
              unloadMuxOut[1] = fifoOut[16][11][w-1];
              unloadMuxOut[2] = fifoOut[17][11][w-1];
              unloadMuxOut[3] = fifoOut[18][11][w-1];
              unloadMuxOut[4] = fifoOut[19][11][w-1];
              unloadMuxOut[5] = fifoOut[20][11][w-1];
              unloadMuxOut[6] = fifoOut[21][11][w-1];
              unloadMuxOut[7] = fifoOut[22][11][w-1];
              unloadMuxOut[8] = fifoOut[23][11][w-1];
              unloadMuxOut[9] = fifoOut[24][11][w-1];
              unloadMuxOut[10] = fifoOut[25][11][w-1];
              unloadMuxOut[11] = fifoOut[0][10][w-1];
              unloadMuxOut[12] = fifoOut[1][10][w-1];
              unloadMuxOut[13] = fifoOut[2][10][w-1];
              unloadMuxOut[14] = fifoOut[3][10][w-1];
              unloadMuxOut[15] = fifoOut[4][10][w-1];
              unloadMuxOut[16] = fifoOut[5][10][w-1];
              unloadMuxOut[17] = fifoOut[6][10][w-1];
              unloadMuxOut[18] = fifoOut[7][10][w-1];
              unloadMuxOut[19] = fifoOut[8][10][w-1];
              unloadMuxOut[20] = fifoOut[9][10][w-1];
              unloadMuxOut[21] = fifoOut[10][10][w-1];
              unloadMuxOut[22] = fifoOut[11][10][w-1];
              unloadMuxOut[23] = fifoOut[12][10][w-1];
              unloadMuxOut[24] = fifoOut[13][10][w-1];
              unloadMuxOut[25] = fifoOut[14][10][w-1];
              unloadMuxOut[26] = fifoOut[15][10][w-1];
              unloadMuxOut[27] = fifoOut[16][10][w-1];
              unloadMuxOut[28] = fifoOut[17][10][w-1];
              unloadMuxOut[29] = fifoOut[18][10][w-1];
              unloadMuxOut[30] = fifoOut[19][10][w-1];
              unloadMuxOut[31] = fifoOut[20][10][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[21][10][w-1];
              unloadMuxOut[1] = fifoOut[22][10][w-1];
              unloadMuxOut[2] = fifoOut[23][10][w-1];
              unloadMuxOut[3] = fifoOut[24][10][w-1];
              unloadMuxOut[4] = fifoOut[25][10][w-1];
              unloadMuxOut[5] = fifoOut[0][9][w-1];
              unloadMuxOut[6] = fifoOut[1][9][w-1];
              unloadMuxOut[7] = fifoOut[2][9][w-1];
              unloadMuxOut[8] = fifoOut[3][9][w-1];
              unloadMuxOut[9] = fifoOut[4][9][w-1];
              unloadMuxOut[10] = fifoOut[5][9][w-1];
              unloadMuxOut[11] = fifoOut[6][9][w-1];
              unloadMuxOut[12] = fifoOut[7][9][w-1];
              unloadMuxOut[13] = fifoOut[8][9][w-1];
              unloadMuxOut[14] = fifoOut[9][9][w-1];
              unloadMuxOut[15] = fifoOut[10][9][w-1];
              unloadMuxOut[16] = fifoOut[11][9][w-1];
              unloadMuxOut[17] = fifoOut[12][9][w-1];
              unloadMuxOut[18] = fifoOut[13][9][w-1];
              unloadMuxOut[19] = fifoOut[14][9][w-1];
              unloadMuxOut[20] = fifoOut[15][9][w-1];
              unloadMuxOut[21] = fifoOut[16][9][w-1];
              unloadMuxOut[22] = fifoOut[17][9][w-1];
              unloadMuxOut[23] = fifoOut[18][9][w-1];
              unloadMuxOut[24] = fifoOut[19][9][w-1];
              unloadMuxOut[25] = fifoOut[20][9][w-1];
              unloadMuxOut[26] = fifoOut[21][9][w-1];
              unloadMuxOut[27] = fifoOut[22][9][w-1];
              unloadMuxOut[28] = fifoOut[23][9][w-1];
              unloadMuxOut[29] = fifoOut[24][9][w-1];
              unloadMuxOut[30] = fifoOut[25][9][w-1];
              unloadMuxOut[31] = fifoOut[0][8][w-1];
       end
       16: begin
              unloadMuxOut[0] = fifoOut[1][8][w-1];
              unloadMuxOut[1] = fifoOut[2][8][w-1];
              unloadMuxOut[2] = fifoOut[3][8][w-1];
              unloadMuxOut[3] = fifoOut[4][8][w-1];
              unloadMuxOut[4] = fifoOut[5][8][w-1];
              unloadMuxOut[5] = fifoOut[6][8][w-1];
              unloadMuxOut[6] = fifoOut[7][8][w-1];
              unloadMuxOut[7] = fifoOut[8][8][w-1];
              unloadMuxOut[8] = fifoOut[9][8][w-1];
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0; 
             end
       end
    endcase //unload case end
         case(rd_address_case)
         0: begin
              muxOutConnector[0] = fifoOut[10][8];
              muxOutConnector[1] = fifoOut[11][8];
              muxOutConnector[2] = fifoOut[12][8];
              muxOutConnector[3] = fifoOut[13][8];
              muxOutConnector[4] = fifoOut[14][8];
              muxOutConnector[5] = fifoOut[15][8];
              muxOutConnector[6] = fifoOut[16][8];
              muxOutConnector[7] = fifoOut[17][8];
              muxOutConnector[8] = fifoOut[18][8];
              muxOutConnector[9] = fifoOut[19][8];
              muxOutConnector[10] = fifoOut[20][8];
              muxOutConnector[11] = fifoOut[21][8];
              muxOutConnector[12] = fifoOut[22][8];
              muxOutConnector[13] = fifoOut[23][8];
              muxOutConnector[14] = fifoOut[24][8];
              muxOutConnector[15] = fifoOut[25][8];
              muxOutConnector[16] = fifoOut[0][7];
              muxOutConnector[17] = fifoOut[1][7];
              muxOutConnector[18] = fifoOut[2][7];
              muxOutConnector[19] = fifoOut[3][7];
              muxOutConnector[20] = fifoOut[4][7];
              muxOutConnector[21] = fifoOut[5][7];
              muxOutConnector[22] = fifoOut[6][7];
              muxOutConnector[23] = fifoOut[7][7];
              muxOutConnector[24] = fifoOut[8][7];
              muxOutConnector[25] = fifoOut[9][7];
              muxOutConnector[26] = fifoOut[41][1];
              muxOutConnector[27] = fifoOut[42][1];
              muxOutConnector[28] = fifoOut[43][1];
              muxOutConnector[29] = fifoOut[44][1];
              muxOutConnector[30] = fifoOut[45][1];
              muxOutConnector[31] = fifoOut[46][1];
              muxOutConnector[32] = fifoOut[47][1];
              muxOutConnector[33] = fifoOut[48][1];
              muxOutConnector[34] = fifoOut[49][1];
              muxOutConnector[35] = fifoOut[50][1];
              muxOutConnector[36] = fifoOut[51][1];
              muxOutConnector[37] = fifoOut[26][0];
              muxOutConnector[38] = fifoOut[27][0];
              muxOutConnector[39] = fifoOut[28][0];
              muxOutConnector[40] = fifoOut[29][0];
              muxOutConnector[41] = fifoOut[30][0];
              muxOutConnector[42] = fifoOut[31][0];
              muxOutConnector[43] = fifoOut[32][0];
              muxOutConnector[44] = fifoOut[33][0];
              muxOutConnector[45] = fifoOut[34][0];
              muxOutConnector[46] = fifoOut[35][0];
              muxOutConnector[47] = fifoOut[36][0];
              muxOutConnector[48] = fifoOut[37][0];
              muxOutConnector[49] = fifoOut[38][0];
              muxOutConnector[50] = fifoOut[39][0];
              muxOutConnector[51] = fifoOut[40][0];
         end
         1: begin
              muxOutConnector[0] = fifoOut[10][7];
              muxOutConnector[1] = fifoOut[11][7];
              muxOutConnector[2] = fifoOut[12][7];
              muxOutConnector[3] = fifoOut[13][7];
              muxOutConnector[4] = fifoOut[14][7];
              muxOutConnector[5] = fifoOut[15][7];
              muxOutConnector[6] = fifoOut[16][7];
              muxOutConnector[7] = fifoOut[17][7];
              muxOutConnector[8] = fifoOut[18][7];
              muxOutConnector[9] = fifoOut[19][7];
              muxOutConnector[10] = fifoOut[20][7];
              muxOutConnector[11] = fifoOut[21][7];
              muxOutConnector[12] = fifoOut[22][7];
              muxOutConnector[13] = fifoOut[23][7];
              muxOutConnector[14] = fifoOut[24][7];
              muxOutConnector[15] = fifoOut[25][7];
              muxOutConnector[16] = fifoOut[0][6];
              muxOutConnector[17] = fifoOut[1][6];
              muxOutConnector[18] = fifoOut[2][6];
              muxOutConnector[19] = fifoOut[3][6];
              muxOutConnector[20] = fifoOut[4][6];
              muxOutConnector[21] = fifoOut[5][6];
              muxOutConnector[22] = fifoOut[6][6];
              muxOutConnector[23] = fifoOut[7][6];
              muxOutConnector[24] = fifoOut[8][6];
              muxOutConnector[25] = fifoOut[9][6];
              muxOutConnector[26] = fifoOut[41][0];
              muxOutConnector[27] = fifoOut[42][0];
              muxOutConnector[28] = fifoOut[23][12];
              muxOutConnector[29] = fifoOut[24][12];
              muxOutConnector[30] = fifoOut[25][12];
              muxOutConnector[31] = fifoOut[0][11];
              muxOutConnector[32] = fifoOut[1][11];
              muxOutConnector[33] = fifoOut[2][11];
              muxOutConnector[34] = fifoOut[3][11];
              muxOutConnector[35] = fifoOut[4][11];
              muxOutConnector[36] = fifoOut[5][11];
              muxOutConnector[37] = fifoOut[6][11];
              muxOutConnector[38] = fifoOut[7][11];
              muxOutConnector[39] = fifoOut[8][11];
              muxOutConnector[40] = fifoOut[9][11];
              muxOutConnector[41] = fifoOut[10][11];
              muxOutConnector[42] = fifoOut[11][11];
              muxOutConnector[43] = fifoOut[12][11];
              muxOutConnector[44] = fifoOut[13][11];
              muxOutConnector[45] = fifoOut[14][11];
              muxOutConnector[46] = fifoOut[15][11];
              muxOutConnector[47] = fifoOut[16][11];
              muxOutConnector[48] = fifoOut[17][11];
              muxOutConnector[49] = fifoOut[18][11];
              muxOutConnector[50] = fifoOut[19][11];
              muxOutConnector[51] = fifoOut[20][11];
         end
         2: begin
              muxOutConnector[0] = fifoOut[10][6];
              muxOutConnector[1] = fifoOut[11][6];
              muxOutConnector[2] = fifoOut[12][6];
              muxOutConnector[3] = fifoOut[13][6];
              muxOutConnector[4] = fifoOut[14][6];
              muxOutConnector[5] = fifoOut[15][6];
              muxOutConnector[6] = fifoOut[16][6];
              muxOutConnector[7] = fifoOut[17][6];
              muxOutConnector[8] = fifoOut[18][6];
              muxOutConnector[9] = fifoOut[19][6];
              muxOutConnector[10] = fifoOut[20][6];
              muxOutConnector[11] = fifoOut[21][6];
              muxOutConnector[12] = fifoOut[22][6];
              muxOutConnector[13] = fifoOut[23][6];
              muxOutConnector[14] = fifoOut[24][6];
              muxOutConnector[15] = fifoOut[25][6];
              muxOutConnector[16] = fifoOut[0][5];
              muxOutConnector[17] = fifoOut[1][5];
              muxOutConnector[18] = fifoOut[2][5];
              muxOutConnector[19] = fifoOut[3][5];
              muxOutConnector[20] = fifoOut[4][5];
              muxOutConnector[21] = fifoOut[5][5];
              muxOutConnector[22] = fifoOut[6][5];
              muxOutConnector[23] = fifoOut[7][5];
              muxOutConnector[24] = fifoOut[8][5];
              muxOutConnector[25] = fifoOut[9][5];
              muxOutConnector[26] = fifoOut[21][11];
              muxOutConnector[27] = fifoOut[22][11];
              muxOutConnector[28] = fifoOut[23][11];
              muxOutConnector[29] = fifoOut[24][11];
              muxOutConnector[30] = fifoOut[25][11];
              muxOutConnector[31] = fifoOut[0][10];
              muxOutConnector[32] = fifoOut[1][10];
              muxOutConnector[33] = fifoOut[2][10];
              muxOutConnector[34] = fifoOut[3][10];
              muxOutConnector[35] = fifoOut[4][10];
              muxOutConnector[36] = fifoOut[5][10];
              muxOutConnector[37] = fifoOut[6][10];
              muxOutConnector[38] = fifoOut[7][10];
              muxOutConnector[39] = fifoOut[8][10];
              muxOutConnector[40] = fifoOut[9][10];
              muxOutConnector[41] = fifoOut[10][10];
              muxOutConnector[42] = fifoOut[11][10];
              muxOutConnector[43] = fifoOut[12][10];
              muxOutConnector[44] = fifoOut[13][10];
              muxOutConnector[45] = fifoOut[14][10];
              muxOutConnector[46] = fifoOut[15][10];
              muxOutConnector[47] = fifoOut[16][10];
              muxOutConnector[48] = fifoOut[17][10];
              muxOutConnector[49] = fifoOut[18][10];
              muxOutConnector[50] = fifoOut[19][10];
              muxOutConnector[51] = fifoOut[20][10];
         end
         3: begin
              muxOutConnector[0] = fifoOut[10][5];
              muxOutConnector[1] = fifoOut[11][5];
              muxOutConnector[2] = fifoOut[12][5];
              muxOutConnector[3] = fifoOut[13][5];
              muxOutConnector[4] = fifoOut[14][5];
              muxOutConnector[5] = fifoOut[15][5];
              muxOutConnector[6] = fifoOut[16][5];
              muxOutConnector[7] = fifoOut[17][5];
              muxOutConnector[8] = fifoOut[18][5];
              muxOutConnector[9] = fifoOut[19][5];
              muxOutConnector[10] = fifoOut[20][5];
              muxOutConnector[11] = fifoOut[21][5];
              muxOutConnector[12] = fifoOut[22][5];
              muxOutConnector[13] = fifoOut[23][5];
              muxOutConnector[14] = fifoOut[24][5];
              muxOutConnector[15] = fifoOut[25][5];
              muxOutConnector[16] = fifoOut[0][4];
              muxOutConnector[17] = fifoOut[1][4];
              muxOutConnector[18] = fifoOut[2][4];
              muxOutConnector[19] = fifoOut[3][4];
              muxOutConnector[20] = fifoOut[4][4];
              muxOutConnector[21] = fifoOut[5][4];
              muxOutConnector[22] = fifoOut[6][4];
              muxOutConnector[23] = fifoOut[7][4];
              muxOutConnector[24] = fifoOut[8][4];
              muxOutConnector[25] = fifoOut[9][4];
              muxOutConnector[26] = fifoOut[21][10];
              muxOutConnector[27] = fifoOut[22][10];
              muxOutConnector[28] = fifoOut[23][10];
              muxOutConnector[29] = fifoOut[24][10];
              muxOutConnector[30] = fifoOut[25][10];
              muxOutConnector[31] = fifoOut[0][9];
              muxOutConnector[32] = fifoOut[1][9];
              muxOutConnector[33] = fifoOut[2][9];
              muxOutConnector[34] = fifoOut[3][9];
              muxOutConnector[35] = fifoOut[4][9];
              muxOutConnector[36] = fifoOut[5][9];
              muxOutConnector[37] = fifoOut[6][9];
              muxOutConnector[38] = fifoOut[7][9];
              muxOutConnector[39] = fifoOut[8][9];
              muxOutConnector[40] = fifoOut[9][9];
              muxOutConnector[41] = fifoOut[10][9];
              muxOutConnector[42] = fifoOut[11][9];
              muxOutConnector[43] = fifoOut[12][9];
              muxOutConnector[44] = fifoOut[13][9];
              muxOutConnector[45] = fifoOut[14][9];
              muxOutConnector[46] = fifoOut[15][9];
              muxOutConnector[47] = fifoOut[16][9];
              muxOutConnector[48] = fifoOut[17][9];
              muxOutConnector[49] = fifoOut[18][9];
              muxOutConnector[50] = fifoOut[19][9];
              muxOutConnector[51] = fifoOut[20][9];
         end
         4: begin
              muxOutConnector[0] = fifoOut[10][4];
              muxOutConnector[1] = fifoOut[11][4];
              muxOutConnector[2] = fifoOut[12][4];
              muxOutConnector[3] = fifoOut[13][4];
              muxOutConnector[4] = fifoOut[14][4];
              muxOutConnector[5] = fifoOut[15][4];
              muxOutConnector[6] = fifoOut[16][4];
              muxOutConnector[7] = fifoOut[17][4];
              muxOutConnector[8] = fifoOut[18][4];
              muxOutConnector[9] = fifoOut[19][4];
              muxOutConnector[10] = fifoOut[20][4];
              muxOutConnector[11] = fifoOut[21][4];
              muxOutConnector[12] = fifoOut[22][4];
              muxOutConnector[13] = fifoOut[23][4];
              muxOutConnector[14] = fifoOut[24][4];
              muxOutConnector[15] = fifoOut[25][4];
              muxOutConnector[16] = fifoOut[0][3];
              muxOutConnector[17] = fifoOut[1][3];
              muxOutConnector[18] = fifoOut[2][3];
              muxOutConnector[19] = fifoOut[3][3];
              muxOutConnector[20] = fifoOut[4][3];
              muxOutConnector[21] = fifoOut[5][3];
              muxOutConnector[22] = fifoOut[6][3];
              muxOutConnector[23] = fifoOut[7][3];
              muxOutConnector[24] = fifoOut[8][3];
              muxOutConnector[25] = fifoOut[9][3];
              muxOutConnector[26] = fifoOut[21][9];
              muxOutConnector[27] = fifoOut[22][9];
              muxOutConnector[28] = fifoOut[23][9];
              muxOutConnector[29] = fifoOut[24][9];
              muxOutConnector[30] = fifoOut[25][9];
              muxOutConnector[31] = fifoOut[0][8];
              muxOutConnector[32] = fifoOut[1][8];
              muxOutConnector[33] = fifoOut[2][8];
              muxOutConnector[34] = fifoOut[3][8];
              muxOutConnector[35] = fifoOut[4][8];
              muxOutConnector[36] = fifoOut[5][8];
              muxOutConnector[37] = fifoOut[6][8];
              muxOutConnector[38] = fifoOut[7][8];
              muxOutConnector[39] = fifoOut[8][8];
              muxOutConnector[40] = fifoOut[9][8];
              muxOutConnector[41] = fifoOut[10][8];
              muxOutConnector[42] = fifoOut[11][8];
              muxOutConnector[43] = fifoOut[12][8];
              muxOutConnector[44] = fifoOut[13][8];
              muxOutConnector[45] = fifoOut[14][8];
              muxOutConnector[46] = fifoOut[15][8];
              muxOutConnector[47] = fifoOut[16][8];
              muxOutConnector[48] = fifoOut[17][8];
              muxOutConnector[49] = fifoOut[18][8];
              muxOutConnector[50] = fifoOut[19][8];
              muxOutConnector[51] = fifoOut[20][8];
         end
         5: begin
              muxOutConnector[0] = fifoOut[10][3];
              muxOutConnector[1] = fifoOut[11][3];
              muxOutConnector[2] = fifoOut[12][3];
              muxOutConnector[3] = fifoOut[13][3];
              muxOutConnector[4] = fifoOut[14][3];
              muxOutConnector[5] = fifoOut[15][3];
              muxOutConnector[6] = fifoOut[16][3];
              muxOutConnector[7] = fifoOut[17][3];
              muxOutConnector[8] = fifoOut[18][3];
              muxOutConnector[9] = fifoOut[19][3];
              muxOutConnector[10] = fifoOut[20][3];
              muxOutConnector[11] = fifoOut[21][3];
              muxOutConnector[12] = fifoOut[22][3];
              muxOutConnector[13] = fifoOut[23][3];
              muxOutConnector[14] = fifoOut[24][3];
              muxOutConnector[15] = fifoOut[25][3];
              muxOutConnector[16] = fifoOut[0][2];
              muxOutConnector[17] = fifoOut[1][2];
              muxOutConnector[18] = fifoOut[2][2];
              muxOutConnector[19] = fifoOut[3][2];
              muxOutConnector[20] = fifoOut[4][2];
              muxOutConnector[21] = fifoOut[5][2];
              muxOutConnector[22] = fifoOut[6][2];
              muxOutConnector[23] = fifoOut[7][2];
              muxOutConnector[24] = fifoOut[8][2];
              muxOutConnector[25] = fifoOut[9][2];
              muxOutConnector[26] = fifoOut[21][8];
              muxOutConnector[27] = fifoOut[22][8];
              muxOutConnector[28] = fifoOut[23][8];
              muxOutConnector[29] = fifoOut[24][8];
              muxOutConnector[30] = fifoOut[25][8];
              muxOutConnector[31] = fifoOut[0][7];
              muxOutConnector[32] = fifoOut[1][7];
              muxOutConnector[33] = fifoOut[2][7];
              muxOutConnector[34] = fifoOut[3][7];
              muxOutConnector[35] = fifoOut[4][7];
              muxOutConnector[36] = fifoOut[5][7];
              muxOutConnector[37] = fifoOut[6][7];
              muxOutConnector[38] = fifoOut[7][7];
              muxOutConnector[39] = fifoOut[8][7];
              muxOutConnector[40] = fifoOut[9][7];
              muxOutConnector[41] = fifoOut[10][7];
              muxOutConnector[42] = fifoOut[11][7];
              muxOutConnector[43] = fifoOut[12][7];
              muxOutConnector[44] = fifoOut[13][7];
              muxOutConnector[45] = fifoOut[14][7];
              muxOutConnector[46] = fifoOut[15][7];
              muxOutConnector[47] = fifoOut[16][7];
              muxOutConnector[48] = fifoOut[17][7];
              muxOutConnector[49] = fifoOut[18][7];
              muxOutConnector[50] = fifoOut[19][7];
              muxOutConnector[51] = fifoOut[20][7];
         end
         6: begin
              muxOutConnector[0] = fifoOut[10][2];
              muxOutConnector[1] = fifoOut[11][2];
              muxOutConnector[2] = fifoOut[12][2];
              muxOutConnector[3] = fifoOut[13][2];
              muxOutConnector[4] = fifoOut[14][2];
              muxOutConnector[5] = fifoOut[15][2];
              muxOutConnector[6] = fifoOut[16][2];
              muxOutConnector[7] = fifoOut[17][2];
              muxOutConnector[8] = fifoOut[18][2];
              muxOutConnector[9] = fifoOut[19][2];
              muxOutConnector[10] = fifoOut[20][2];
              muxOutConnector[11] = fifoOut[21][2];
              muxOutConnector[12] = fifoOut[22][2];
              muxOutConnector[13] = fifoOut[23][2];
              muxOutConnector[14] = fifoOut[24][2];
              muxOutConnector[15] = fifoOut[25][2];
              muxOutConnector[16] = fifoOut[0][1];
              muxOutConnector[17] = fifoOut[1][1];
              muxOutConnector[18] = fifoOut[2][1];
              muxOutConnector[19] = fifoOut[3][1];
              muxOutConnector[20] = fifoOut[4][1];
              muxOutConnector[21] = fifoOut[5][1];
              muxOutConnector[22] = fifoOut[6][1];
              muxOutConnector[23] = fifoOut[7][1];
              muxOutConnector[24] = fifoOut[8][1];
              muxOutConnector[25] = fifoOut[9][1];
              muxOutConnector[26] = fifoOut[21][7];
              muxOutConnector[27] = fifoOut[22][7];
              muxOutConnector[28] = fifoOut[23][7];
              muxOutConnector[29] = fifoOut[24][7];
              muxOutConnector[30] = fifoOut[25][7];
              muxOutConnector[31] = fifoOut[0][6];
              muxOutConnector[32] = fifoOut[1][6];
              muxOutConnector[33] = fifoOut[2][6];
              muxOutConnector[34] = fifoOut[3][6];
              muxOutConnector[35] = fifoOut[4][6];
              muxOutConnector[36] = fifoOut[5][6];
              muxOutConnector[37] = fifoOut[6][6];
              muxOutConnector[38] = fifoOut[7][6];
              muxOutConnector[39] = fifoOut[8][6];
              muxOutConnector[40] = fifoOut[9][6];
              muxOutConnector[41] = fifoOut[10][6];
              muxOutConnector[42] = fifoOut[11][6];
              muxOutConnector[43] = fifoOut[12][6];
              muxOutConnector[44] = fifoOut[13][6];
              muxOutConnector[45] = fifoOut[14][6];
              muxOutConnector[46] = fifoOut[15][6];
              muxOutConnector[47] = fifoOut[16][6];
              muxOutConnector[48] = fifoOut[17][6];
              muxOutConnector[49] = fifoOut[18][6];
              muxOutConnector[50] = fifoOut[19][6];
              muxOutConnector[51] = fifoOut[20][6];
         end
         7: begin
              muxOutConnector[0] = fifoOut[10][1];
              muxOutConnector[1] = fifoOut[11][1];
              muxOutConnector[2] = fifoOut[12][1];
              muxOutConnector[3] = fifoOut[13][1];
              muxOutConnector[4] = fifoOut[14][1];
              muxOutConnector[5] = fifoOut[15][1];
              muxOutConnector[6] = fifoOut[16][1];
              muxOutConnector[7] = fifoOut[17][1];
              muxOutConnector[8] = fifoOut[18][1];
              muxOutConnector[9] = fifoOut[19][1];
              muxOutConnector[10] = fifoOut[20][1];
              muxOutConnector[11] = fifoOut[21][1];
              muxOutConnector[12] = fifoOut[22][1];
              muxOutConnector[13] = fifoOut[23][1];
              muxOutConnector[14] = fifoOut[24][1];
              muxOutConnector[15] = fifoOut[25][1];
              muxOutConnector[16] = fifoOut[0][0];
              muxOutConnector[17] = fifoOut[1][0];
              muxOutConnector[18] = fifoOut[2][0];
              muxOutConnector[19] = fifoOut[3][0];
              muxOutConnector[20] = fifoOut[4][0];
              muxOutConnector[21] = fifoOut[5][0];
              muxOutConnector[22] = fifoOut[6][0];
              muxOutConnector[23] = fifoOut[7][0];
              muxOutConnector[24] = fifoOut[8][0];
              muxOutConnector[25] = fifoOut[9][0];
              muxOutConnector[26] = fifoOut[21][6];
              muxOutConnector[27] = fifoOut[22][6];
              muxOutConnector[28] = fifoOut[23][6];
              muxOutConnector[29] = fifoOut[24][6];
              muxOutConnector[30] = fifoOut[25][6];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = fifoOut[12][5];
              muxOutConnector[44] = fifoOut[13][5];
              muxOutConnector[45] = fifoOut[14][5];
              muxOutConnector[46] = fifoOut[15][5];
              muxOutConnector[47] = fifoOut[16][5];
              muxOutConnector[48] = fifoOut[17][5];
              muxOutConnector[49] = fifoOut[18][5];
              muxOutConnector[50] = fifoOut[19][5];
              muxOutConnector[51] = fifoOut[20][5];
         end
         8: begin
              muxOutConnector[0] = fifoOut[10][0];
              muxOutConnector[1] = fifoOut[11][0];
              muxOutConnector[2] = fifoOut[12][0];
              muxOutConnector[3] = fifoOut[13][0];
              muxOutConnector[4] = fifoOut[14][0];
              muxOutConnector[5] = fifoOut[15][0];
              muxOutConnector[6] = fifoOut[16][0];
              muxOutConnector[7] = fifoOut[46][8];
              muxOutConnector[8] = fifoOut[47][8];
              muxOutConnector[9] = fifoOut[48][8];
              muxOutConnector[10] = fifoOut[49][8];
              muxOutConnector[11] = fifoOut[50][8];
              muxOutConnector[12] = fifoOut[51][8];
              muxOutConnector[13] = fifoOut[26][7];
              muxOutConnector[14] = fifoOut[27][7];
              muxOutConnector[15] = fifoOut[28][7];
              muxOutConnector[16] = fifoOut[29][7];
              muxOutConnector[17] = fifoOut[30][7];
              muxOutConnector[18] = fifoOut[31][7];
              muxOutConnector[19] = fifoOut[32][7];
              muxOutConnector[20] = fifoOut[33][7];
              muxOutConnector[21] = fifoOut[34][7];
              muxOutConnector[22] = fifoOut[35][7];
              muxOutConnector[23] = fifoOut[36][7];
              muxOutConnector[24] = fifoOut[37][7];
              muxOutConnector[25] = fifoOut[38][7];
              muxOutConnector[26] = fifoOut[21][5];
              muxOutConnector[27] = fifoOut[22][5];
              muxOutConnector[28] = fifoOut[23][5];
              muxOutConnector[29] = fifoOut[24][5];
              muxOutConnector[30] = fifoOut[25][5];
              muxOutConnector[31] = fifoOut[0][4];
              muxOutConnector[32] = fifoOut[1][4];
              muxOutConnector[33] = fifoOut[2][4];
              muxOutConnector[34] = fifoOut[3][4];
              muxOutConnector[35] = fifoOut[4][4];
              muxOutConnector[36] = fifoOut[5][4];
              muxOutConnector[37] = fifoOut[6][4];
              muxOutConnector[38] = fifoOut[7][4];
              muxOutConnector[39] = fifoOut[8][4];
              muxOutConnector[40] = fifoOut[9][4];
              muxOutConnector[41] = fifoOut[10][4];
              muxOutConnector[42] = fifoOut[11][4];
              muxOutConnector[43] = fifoOut[12][4];
              muxOutConnector[44] = fifoOut[13][4];
              muxOutConnector[45] = fifoOut[14][4];
              muxOutConnector[46] = fifoOut[15][4];
              muxOutConnector[47] = fifoOut[16][4];
              muxOutConnector[48] = fifoOut[17][4];
              muxOutConnector[49] = fifoOut[18][4];
              muxOutConnector[50] = fifoOut[19][4];
              muxOutConnector[51] = fifoOut[20][4];
         end
         9: begin
              muxOutConnector[0] = fifoOut[39][7];
              muxOutConnector[1] = fifoOut[40][7];
              muxOutConnector[2] = fifoOut[41][7];
              muxOutConnector[3] = fifoOut[42][7];
              muxOutConnector[4] = fifoOut[43][7];
              muxOutConnector[5] = fifoOut[44][7];
              muxOutConnector[6] = fifoOut[45][7];
              muxOutConnector[7] = fifoOut[46][7];
              muxOutConnector[8] = fifoOut[47][7];
              muxOutConnector[9] = fifoOut[48][7];
              muxOutConnector[10] = fifoOut[49][7];
              muxOutConnector[11] = fifoOut[50][7];
              muxOutConnector[12] = fifoOut[51][7];
              muxOutConnector[13] = fifoOut[26][6];
              muxOutConnector[14] = fifoOut[27][6];
              muxOutConnector[15] = fifoOut[28][6];
              muxOutConnector[16] = fifoOut[29][6];
              muxOutConnector[17] = fifoOut[30][6];
              muxOutConnector[18] = fifoOut[31][6];
              muxOutConnector[19] = fifoOut[32][6];
              muxOutConnector[20] = fifoOut[33][6];
              muxOutConnector[21] = fifoOut[34][6];
              muxOutConnector[22] = fifoOut[35][6];
              muxOutConnector[23] = fifoOut[36][6];
              muxOutConnector[24] = fifoOut[37][6];
              muxOutConnector[25] = fifoOut[38][6];
              muxOutConnector[26] = fifoOut[21][4];
              muxOutConnector[27] = fifoOut[22][4];
              muxOutConnector[28] = fifoOut[23][4];
              muxOutConnector[29] = fifoOut[24][4];
              muxOutConnector[30] = fifoOut[25][4];
              muxOutConnector[31] = fifoOut[0][3];
              muxOutConnector[32] = fifoOut[1][3];
              muxOutConnector[33] = fifoOut[2][3];
              muxOutConnector[34] = fifoOut[3][3];
              muxOutConnector[35] = fifoOut[4][3];
              muxOutConnector[36] = fifoOut[5][3];
              muxOutConnector[37] = fifoOut[6][3];
              muxOutConnector[38] = fifoOut[7][3];
              muxOutConnector[39] = fifoOut[8][3];
              muxOutConnector[40] = fifoOut[9][3];
              muxOutConnector[41] = fifoOut[10][3];
              muxOutConnector[42] = fifoOut[11][3];
              muxOutConnector[43] = fifoOut[12][3];
              muxOutConnector[44] = fifoOut[13][3];
              muxOutConnector[45] = fifoOut[14][3];
              muxOutConnector[46] = fifoOut[15][3];
              muxOutConnector[47] = fifoOut[16][3];
              muxOutConnector[48] = fifoOut[17][3];
              muxOutConnector[49] = fifoOut[18][3];
              muxOutConnector[50] = fifoOut[19][3];
              muxOutConnector[51] = fifoOut[20][3];
         end
         10: begin
              muxOutConnector[0] = fifoOut[39][6];
              muxOutConnector[1] = fifoOut[40][6];
              muxOutConnector[2] = fifoOut[41][6];
              muxOutConnector[3] = fifoOut[42][6];
              muxOutConnector[4] = fifoOut[43][6];
              muxOutConnector[5] = fifoOut[44][6];
              muxOutConnector[6] = fifoOut[45][6];
              muxOutConnector[7] = fifoOut[46][6];
              muxOutConnector[8] = fifoOut[47][6];
              muxOutConnector[9] = fifoOut[48][6];
              muxOutConnector[10] = fifoOut[49][6];
              muxOutConnector[11] = fifoOut[50][6];
              muxOutConnector[12] = fifoOut[51][6];
              muxOutConnector[13] = fifoOut[26][5];
              muxOutConnector[14] = fifoOut[27][5];
              muxOutConnector[15] = fifoOut[28][5];
              muxOutConnector[16] = fifoOut[29][5];
              muxOutConnector[17] = fifoOut[30][5];
              muxOutConnector[18] = fifoOut[31][5];
              muxOutConnector[19] = fifoOut[32][5];
              muxOutConnector[20] = fifoOut[33][5];
              muxOutConnector[21] = fifoOut[34][5];
              muxOutConnector[22] = fifoOut[35][5];
              muxOutConnector[23] = fifoOut[36][5];
              muxOutConnector[24] = fifoOut[37][5];
              muxOutConnector[25] = fifoOut[38][5];
              muxOutConnector[26] = fifoOut[21][3];
              muxOutConnector[27] = fifoOut[22][3];
              muxOutConnector[28] = fifoOut[23][3];
              muxOutConnector[29] = fifoOut[24][3];
              muxOutConnector[30] = fifoOut[25][3];
              muxOutConnector[31] = fifoOut[0][2];
              muxOutConnector[32] = fifoOut[1][2];
              muxOutConnector[33] = fifoOut[2][2];
              muxOutConnector[34] = fifoOut[3][2];
              muxOutConnector[35] = fifoOut[4][2];
              muxOutConnector[36] = fifoOut[5][2];
              muxOutConnector[37] = fifoOut[6][2];
              muxOutConnector[38] = fifoOut[7][2];
              muxOutConnector[39] = fifoOut[8][2];
              muxOutConnector[40] = fifoOut[9][2];
              muxOutConnector[41] = fifoOut[10][2];
              muxOutConnector[42] = fifoOut[11][2];
              muxOutConnector[43] = fifoOut[12][2];
              muxOutConnector[44] = fifoOut[13][2];
              muxOutConnector[45] = fifoOut[14][2];
              muxOutConnector[46] = fifoOut[15][2];
              muxOutConnector[47] = fifoOut[16][2];
              muxOutConnector[48] = fifoOut[17][2];
              muxOutConnector[49] = fifoOut[18][2];
              muxOutConnector[50] = fifoOut[19][2];
              muxOutConnector[51] = fifoOut[20][2];
         end
         11: begin
              muxOutConnector[0] = fifoOut[39][5];
              muxOutConnector[1] = fifoOut[40][5];
              muxOutConnector[2] = fifoOut[41][5];
              muxOutConnector[3] = fifoOut[42][5];
              muxOutConnector[4] = fifoOut[43][5];
              muxOutConnector[5] = fifoOut[44][5];
              muxOutConnector[6] = fifoOut[45][5];
              muxOutConnector[7] = fifoOut[46][5];
              muxOutConnector[8] = fifoOut[47][5];
              muxOutConnector[9] = fifoOut[48][5];
              muxOutConnector[10] = fifoOut[49][5];
              muxOutConnector[11] = fifoOut[50][5];
              muxOutConnector[12] = fifoOut[51][5];
              muxOutConnector[13] = fifoOut[26][4];
              muxOutConnector[14] = fifoOut[27][4];
              muxOutConnector[15] = fifoOut[28][4];
              muxOutConnector[16] = fifoOut[29][4];
              muxOutConnector[17] = fifoOut[30][4];
              muxOutConnector[18] = fifoOut[31][4];
              muxOutConnector[19] = fifoOut[32][4];
              muxOutConnector[20] = fifoOut[33][4];
              muxOutConnector[21] = fifoOut[34][4];
              muxOutConnector[22] = fifoOut[35][4];
              muxOutConnector[23] = fifoOut[36][4];
              muxOutConnector[24] = fifoOut[37][4];
              muxOutConnector[25] = fifoOut[38][4];
              muxOutConnector[26] = fifoOut[21][2];
              muxOutConnector[27] = fifoOut[22][2];
              muxOutConnector[28] = fifoOut[23][2];
              muxOutConnector[29] = fifoOut[24][2];
              muxOutConnector[30] = fifoOut[25][2];
              muxOutConnector[31] = fifoOut[0][1];
              muxOutConnector[32] = fifoOut[1][1];
              muxOutConnector[33] = fifoOut[2][1];
              muxOutConnector[34] = fifoOut[3][1];
              muxOutConnector[35] = fifoOut[4][1];
              muxOutConnector[36] = fifoOut[5][1];
              muxOutConnector[37] = fifoOut[6][1];
              muxOutConnector[38] = fifoOut[7][1];
              muxOutConnector[39] = fifoOut[8][1];
              muxOutConnector[40] = fifoOut[9][1];
              muxOutConnector[41] = fifoOut[10][1];
              muxOutConnector[42] = fifoOut[11][1];
              muxOutConnector[43] = fifoOut[12][1];
              muxOutConnector[44] = fifoOut[13][1];
              muxOutConnector[45] = fifoOut[14][1];
              muxOutConnector[46] = fifoOut[15][1];
              muxOutConnector[47] = fifoOut[16][1];
              muxOutConnector[48] = fifoOut[17][1];
              muxOutConnector[49] = fifoOut[18][1];
              muxOutConnector[50] = fifoOut[19][1];
              muxOutConnector[51] = fifoOut[20][1];
         end
         12: begin
              muxOutConnector[0] = fifoOut[39][4];
              muxOutConnector[1] = fifoOut[40][4];
              muxOutConnector[2] = fifoOut[41][4];
              muxOutConnector[3] = fifoOut[42][4];
              muxOutConnector[4] = fifoOut[43][4];
              muxOutConnector[5] = fifoOut[44][4];
              muxOutConnector[6] = fifoOut[45][4];
              muxOutConnector[7] = fifoOut[46][4];
              muxOutConnector[8] = fifoOut[47][4];
              muxOutConnector[9] = fifoOut[48][4];
              muxOutConnector[10] = fifoOut[49][4];
              muxOutConnector[11] = fifoOut[50][4];
              muxOutConnector[12] = fifoOut[51][4];
              muxOutConnector[13] = fifoOut[26][3];
              muxOutConnector[14] = fifoOut[27][3];
              muxOutConnector[15] = fifoOut[28][3];
              muxOutConnector[16] = fifoOut[29][3];
              muxOutConnector[17] = fifoOut[30][3];
              muxOutConnector[18] = fifoOut[31][3];
              muxOutConnector[19] = fifoOut[32][3];
              muxOutConnector[20] = fifoOut[33][3];
              muxOutConnector[21] = fifoOut[34][3];
              muxOutConnector[22] = fifoOut[35][3];
              muxOutConnector[23] = fifoOut[36][3];
              muxOutConnector[24] = fifoOut[37][3];
              muxOutConnector[25] = fifoOut[38][3];
              muxOutConnector[26] = fifoOut[21][1];
              muxOutConnector[27] = fifoOut[22][1];
              muxOutConnector[28] = fifoOut[23][1];
              muxOutConnector[29] = fifoOut[24][1];
              muxOutConnector[30] = fifoOut[25][1];
              muxOutConnector[31] = fifoOut[0][0];
              muxOutConnector[32] = fifoOut[1][0];
              muxOutConnector[33] = fifoOut[2][0];
              muxOutConnector[34] = fifoOut[3][0];
              muxOutConnector[35] = fifoOut[4][0];
              muxOutConnector[36] = fifoOut[5][0];
              muxOutConnector[37] = fifoOut[6][0];
              muxOutConnector[38] = fifoOut[7][0];
              muxOutConnector[39] = fifoOut[8][0];
              muxOutConnector[40] = fifoOut[9][0];
              muxOutConnector[41] = fifoOut[10][0];
              muxOutConnector[42] = fifoOut[11][0];
              muxOutConnector[43] = fifoOut[12][0];
              muxOutConnector[44] = fifoOut[13][0];
              muxOutConnector[45] = fifoOut[14][0];
              muxOutConnector[46] = fifoOut[15][0];
              muxOutConnector[47] = fifoOut[16][0];
              muxOutConnector[48] = fifoOut[46][8];
              muxOutConnector[49] = fifoOut[47][8];
              muxOutConnector[50] = fifoOut[48][8];
              muxOutConnector[51] = fifoOut[49][8];
         end
         13: begin
              muxOutConnector[0] = fifoOut[39][3];
              muxOutConnector[1] = fifoOut[40][3];
              muxOutConnector[2] = fifoOut[41][3];
              muxOutConnector[3] = fifoOut[42][3];
              muxOutConnector[4] = fifoOut[43][3];
              muxOutConnector[5] = fifoOut[44][3];
              muxOutConnector[6] = fifoOut[45][3];
              muxOutConnector[7] = fifoOut[46][3];
              muxOutConnector[8] = fifoOut[47][3];
              muxOutConnector[9] = fifoOut[48][3];
              muxOutConnector[10] = fifoOut[49][3];
              muxOutConnector[11] = fifoOut[50][3];
              muxOutConnector[12] = fifoOut[51][3];
              muxOutConnector[13] = fifoOut[26][2];
              muxOutConnector[14] = fifoOut[27][2];
              muxOutConnector[15] = fifoOut[28][2];
              muxOutConnector[16] = fifoOut[29][2];
              muxOutConnector[17] = fifoOut[30][2];
              muxOutConnector[18] = fifoOut[31][2];
              muxOutConnector[19] = fifoOut[32][2];
              muxOutConnector[20] = fifoOut[33][2];
              muxOutConnector[21] = fifoOut[34][2];
              muxOutConnector[22] = fifoOut[35][2];
              muxOutConnector[23] = fifoOut[36][2];
              muxOutConnector[24] = fifoOut[37][2];
              muxOutConnector[25] = fifoOut[38][2];
              muxOutConnector[26] = fifoOut[50][8];
              muxOutConnector[27] = fifoOut[51][8];
              muxOutConnector[28] = fifoOut[26][7];
              muxOutConnector[29] = fifoOut[27][7];
              muxOutConnector[30] = fifoOut[28][7];
              muxOutConnector[31] = fifoOut[29][7];
              muxOutConnector[32] = fifoOut[30][7];
              muxOutConnector[33] = fifoOut[31][7];
              muxOutConnector[34] = fifoOut[32][7];
              muxOutConnector[35] = fifoOut[33][7];
              muxOutConnector[36] = fifoOut[34][7];
              muxOutConnector[37] = fifoOut[35][7];
              muxOutConnector[38] = fifoOut[36][7];
              muxOutConnector[39] = fifoOut[37][7];
              muxOutConnector[40] = fifoOut[38][7];
              muxOutConnector[41] = fifoOut[39][7];
              muxOutConnector[42] = fifoOut[40][7];
              muxOutConnector[43] = fifoOut[41][7];
              muxOutConnector[44] = fifoOut[42][7];
              muxOutConnector[45] = fifoOut[43][7];
              muxOutConnector[46] = fifoOut[44][7];
              muxOutConnector[47] = fifoOut[45][7];
              muxOutConnector[48] = fifoOut[46][7];
              muxOutConnector[49] = fifoOut[47][7];
              muxOutConnector[50] = fifoOut[48][7];
              muxOutConnector[51] = fifoOut[49][7];
         end
         14: begin
              muxOutConnector[0] = fifoOut[39][2];
              muxOutConnector[1] = fifoOut[40][2];
              muxOutConnector[2] = fifoOut[41][2];
              muxOutConnector[3] = fifoOut[42][2];
              muxOutConnector[4] = fifoOut[43][2];
              muxOutConnector[5] = fifoOut[44][2];
              muxOutConnector[6] = fifoOut[45][2];
              muxOutConnector[7] = fifoOut[46][2];
              muxOutConnector[8] = fifoOut[47][2];
              muxOutConnector[9] = fifoOut[48][2];
              muxOutConnector[10] = fifoOut[49][2];
              muxOutConnector[11] = fifoOut[50][2];
              muxOutConnector[12] = fifoOut[51][2];
              muxOutConnector[13] = fifoOut[26][1];
              muxOutConnector[14] = fifoOut[27][1];
              muxOutConnector[15] = fifoOut[28][1];
              muxOutConnector[16] = fifoOut[29][1];
              muxOutConnector[17] = fifoOut[30][1];
              muxOutConnector[18] = fifoOut[31][1];
              muxOutConnector[19] = fifoOut[32][1];
              muxOutConnector[20] = fifoOut[33][1];
              muxOutConnector[21] = fifoOut[34][1];
              muxOutConnector[22] = fifoOut[35][1];
              muxOutConnector[23] = fifoOut[36][1];
              muxOutConnector[24] = fifoOut[37][1];
              muxOutConnector[25] = fifoOut[38][1];
              muxOutConnector[26] = fifoOut[50][7];
              muxOutConnector[27] = fifoOut[51][7];
              muxOutConnector[28] = fifoOut[26][6];
              muxOutConnector[29] = fifoOut[27][6];
              muxOutConnector[30] = fifoOut[28][6];
              muxOutConnector[31] = fifoOut[29][6];
              muxOutConnector[32] = fifoOut[30][6];
              muxOutConnector[33] = fifoOut[31][6];
              muxOutConnector[34] = fifoOut[32][6];
              muxOutConnector[35] = fifoOut[33][6];
              muxOutConnector[36] = fifoOut[34][6];
              muxOutConnector[37] = fifoOut[35][6];
              muxOutConnector[38] = fifoOut[36][6];
              muxOutConnector[39] = fifoOut[37][6];
              muxOutConnector[40] = fifoOut[38][6];
              muxOutConnector[41] = fifoOut[39][6];
              muxOutConnector[42] = fifoOut[40][6];
              muxOutConnector[43] = fifoOut[41][6];
              muxOutConnector[44] = fifoOut[42][6];
              muxOutConnector[45] = fifoOut[43][6];
              muxOutConnector[46] = fifoOut[44][6];
              muxOutConnector[47] = fifoOut[45][6];
              muxOutConnector[48] = fifoOut[46][6];
              muxOutConnector[49] = fifoOut[47][6];
              muxOutConnector[50] = fifoOut[48][6];
              muxOutConnector[51] = fifoOut[49][6];
         end
         15: begin
              muxOutConnector[0] = fifoOut[39][1];
              muxOutConnector[1] = fifoOut[40][1];
              muxOutConnector[2] = fifoOut[41][1];
              muxOutConnector[3] = fifoOut[42][1];
              muxOutConnector[4] = fifoOut[43][1];
              muxOutConnector[5] = fifoOut[44][1];
              muxOutConnector[6] = fifoOut[45][1];
              muxOutConnector[7] = fifoOut[46][1];
              muxOutConnector[8] = fifoOut[47][1];
              muxOutConnector[9] = fifoOut[48][1];
              muxOutConnector[10] = fifoOut[49][1];
              muxOutConnector[11] = fifoOut[50][1];
              muxOutConnector[12] = fifoOut[51][1];
              muxOutConnector[13] = fifoOut[26][0];
              muxOutConnector[14] = fifoOut[27][0];
              muxOutConnector[15] = fifoOut[28][0];
              muxOutConnector[16] = fifoOut[29][0];
              muxOutConnector[17] = fifoOut[30][0];
              muxOutConnector[18] = fifoOut[31][0];
              muxOutConnector[19] = fifoOut[32][0];
              muxOutConnector[20] = fifoOut[33][0];
              muxOutConnector[21] = fifoOut[34][0];
              muxOutConnector[22] = fifoOut[35][0];
              muxOutConnector[23] = fifoOut[36][0];
              muxOutConnector[24] = fifoOut[37][0];
              muxOutConnector[25] = fifoOut[38][0];
              muxOutConnector[26] = fifoOut[50][6];
              muxOutConnector[27] = fifoOut[51][6];
              muxOutConnector[28] = fifoOut[26][5];
              muxOutConnector[29] = fifoOut[27][5];
              muxOutConnector[30] = fifoOut[28][5];
              muxOutConnector[31] = fifoOut[29][5];
              muxOutConnector[32] = fifoOut[30][5];
              muxOutConnector[33] = fifoOut[31][5];
              muxOutConnector[34] = fifoOut[32][5];
              muxOutConnector[35] = fifoOut[33][5];
              muxOutConnector[36] = fifoOut[34][5];
              muxOutConnector[37] = fifoOut[35][5];
              muxOutConnector[38] = fifoOut[36][5];
              muxOutConnector[39] = fifoOut[37][5];
              muxOutConnector[40] = fifoOut[38][5];
              muxOutConnector[41] = fifoOut[39][5];
              muxOutConnector[42] = fifoOut[40][5];
              muxOutConnector[43] = fifoOut[41][5];
              muxOutConnector[44] = fifoOut[42][5];
              muxOutConnector[45] = fifoOut[43][5];
              muxOutConnector[46] = fifoOut[44][5];
              muxOutConnector[47] = fifoOut[45][5];
              muxOutConnector[48] = fifoOut[46][5];
              muxOutConnector[49] = fifoOut[47][5];
              muxOutConnector[50] = fifoOut[48][5];
              muxOutConnector[51] = fifoOut[49][5];
         end
         16: begin
              muxOutConnector[0] = fifoOut[39][0];
              muxOutConnector[1] = fifoOut[40][0];
              muxOutConnector[2] = fifoOut[41][0];
              muxOutConnector[3] = fifoOut[42][0];
              muxOutConnector[4] = fifoOut[23][12];
              muxOutConnector[5] = fifoOut[24][12];
              muxOutConnector[6] = fifoOut[25][12];
              muxOutConnector[7] = fifoOut[0][11];
              muxOutConnector[8] = fifoOut[1][11];
              muxOutConnector[9] = fifoOut[2][11];
              muxOutConnector[10] = fifoOut[3][11];
              muxOutConnector[11] = fifoOut[4][11];
              muxOutConnector[12] = fifoOut[5][11];
              muxOutConnector[13] = fifoOut[6][11];
              muxOutConnector[14] = fifoOut[7][11];
              muxOutConnector[15] = fifoOut[8][11];
              muxOutConnector[16] = fifoOut[9][11];
              muxOutConnector[17] = fifoOut[10][11];
              muxOutConnector[18] = fifoOut[11][11];
              muxOutConnector[19] = fifoOut[12][11];
              muxOutConnector[20] = fifoOut[13][11];
              muxOutConnector[21] = fifoOut[14][11];
              muxOutConnector[22] = fifoOut[15][11];
              muxOutConnector[23] = fifoOut[16][11];
              muxOutConnector[24] = fifoOut[17][11];
              muxOutConnector[25] = fifoOut[18][11];
              muxOutConnector[26] = fifoOut[50][5];
              muxOutConnector[27] = fifoOut[51][5];
              muxOutConnector[28] = fifoOut[26][4];
              muxOutConnector[29] = fifoOut[27][4];
              muxOutConnector[30] = fifoOut[28][4];
              muxOutConnector[31] = fifoOut[29][4];
              muxOutConnector[32] = fifoOut[30][4];
              muxOutConnector[33] = fifoOut[31][4];
              muxOutConnector[34] = fifoOut[32][4];
              muxOutConnector[35] = fifoOut[33][4];
              muxOutConnector[36] = fifoOut[34][4];
              muxOutConnector[37] = fifoOut[35][4];
              muxOutConnector[38] = fifoOut[36][4];
              muxOutConnector[39] = fifoOut[37][4];
              muxOutConnector[40] = fifoOut[38][4];
              muxOutConnector[41] = fifoOut[39][4];
              muxOutConnector[42] = fifoOut[40][4];
              muxOutConnector[43] = fifoOut[41][4];
              muxOutConnector[44] = fifoOut[42][4];
              muxOutConnector[45] = fifoOut[43][4];
              muxOutConnector[46] = fifoOut[44][4];
              muxOutConnector[47] = fifoOut[45][4];
              muxOutConnector[48] = fifoOut[46][4];
              muxOutConnector[49] = fifoOut[47][4];
              muxOutConnector[50] = fifoOut[48][4];
              muxOutConnector[51] = fifoOut[49][4];
         end
         17: begin
              muxOutConnector[0] = fifoOut[19][11];
              muxOutConnector[1] = fifoOut[20][11];
              muxOutConnector[2] = fifoOut[21][11];
              muxOutConnector[3] = fifoOut[22][11];
              muxOutConnector[4] = fifoOut[23][11];
              muxOutConnector[5] = fifoOut[24][11];
              muxOutConnector[6] = fifoOut[25][11];
              muxOutConnector[7] = fifoOut[0][10];
              muxOutConnector[8] = fifoOut[1][10];
              muxOutConnector[9] = fifoOut[2][10];
              muxOutConnector[10] = fifoOut[3][10];
              muxOutConnector[11] = fifoOut[4][10];
              muxOutConnector[12] = fifoOut[5][10];
              muxOutConnector[13] = fifoOut[6][10];
              muxOutConnector[14] = fifoOut[7][10];
              muxOutConnector[15] = fifoOut[8][10];
              muxOutConnector[16] = fifoOut[9][10];
              muxOutConnector[17] = fifoOut[10][10];
              muxOutConnector[18] = fifoOut[11][10];
              muxOutConnector[19] = fifoOut[12][10];
              muxOutConnector[20] = fifoOut[13][10];
              muxOutConnector[21] = fifoOut[14][10];
              muxOutConnector[22] = fifoOut[15][10];
              muxOutConnector[23] = fifoOut[16][10];
              muxOutConnector[24] = fifoOut[17][10];
              muxOutConnector[25] = fifoOut[18][10];
              muxOutConnector[26] = fifoOut[50][4];
              muxOutConnector[27] = fifoOut[51][4];
              muxOutConnector[28] = fifoOut[26][3];
              muxOutConnector[29] = fifoOut[27][3];
              muxOutConnector[30] = fifoOut[28][3];
              muxOutConnector[31] = fifoOut[29][3];
              muxOutConnector[32] = fifoOut[30][3];
              muxOutConnector[33] = fifoOut[31][3];
              muxOutConnector[34] = fifoOut[32][3];
              muxOutConnector[35] = fifoOut[33][3];
              muxOutConnector[36] = fifoOut[34][3];
              muxOutConnector[37] = fifoOut[35][3];
              muxOutConnector[38] = fifoOut[36][3];
              muxOutConnector[39] = fifoOut[37][3];
              muxOutConnector[40] = fifoOut[38][3];
              muxOutConnector[41] = fifoOut[39][3];
              muxOutConnector[42] = fifoOut[40][3];
              muxOutConnector[43] = fifoOut[41][3];
              muxOutConnector[44] = fifoOut[42][3];
              muxOutConnector[45] = fifoOut[43][3];
              muxOutConnector[46] = fifoOut[44][3];
              muxOutConnector[47] = fifoOut[45][3];
              muxOutConnector[48] = fifoOut[46][3];
              muxOutConnector[49] = fifoOut[47][3];
              muxOutConnector[50] = fifoOut[48][3];
              muxOutConnector[51] = fifoOut[49][3];
         end
         18: begin
              muxOutConnector[0] = fifoOut[19][10];
              muxOutConnector[1] = fifoOut[20][10];
              muxOutConnector[2] = fifoOut[21][10];
              muxOutConnector[3] = fifoOut[22][10];
              muxOutConnector[4] = fifoOut[23][10];
              muxOutConnector[5] = fifoOut[24][10];
              muxOutConnector[6] = fifoOut[25][10];
              muxOutConnector[7] = fifoOut[0][9];
              muxOutConnector[8] = fifoOut[1][9];
              muxOutConnector[9] = fifoOut[2][9];
              muxOutConnector[10] = fifoOut[3][9];
              muxOutConnector[11] = fifoOut[4][9];
              muxOutConnector[12] = fifoOut[5][9];
              muxOutConnector[13] = fifoOut[6][9];
              muxOutConnector[14] = fifoOut[7][9];
              muxOutConnector[15] = fifoOut[8][9];
              muxOutConnector[16] = fifoOut[9][9];
              muxOutConnector[17] = fifoOut[10][9];
              muxOutConnector[18] = fifoOut[11][9];
              muxOutConnector[19] = fifoOut[12][9];
              muxOutConnector[20] = fifoOut[13][9];
              muxOutConnector[21] = fifoOut[14][9];
              muxOutConnector[22] = fifoOut[15][9];
              muxOutConnector[23] = fifoOut[16][9];
              muxOutConnector[24] = fifoOut[17][9];
              muxOutConnector[25] = fifoOut[18][9];
              muxOutConnector[26] = fifoOut[50][3];
              muxOutConnector[27] = fifoOut[51][3];
              muxOutConnector[28] = fifoOut[26][2];
              muxOutConnector[29] = fifoOut[27][2];
              muxOutConnector[30] = fifoOut[28][2];
              muxOutConnector[31] = fifoOut[29][2];
              muxOutConnector[32] = fifoOut[30][2];
              muxOutConnector[33] = fifoOut[31][2];
              muxOutConnector[34] = fifoOut[32][2];
              muxOutConnector[35] = fifoOut[33][2];
              muxOutConnector[36] = fifoOut[34][2];
              muxOutConnector[37] = fifoOut[35][2];
              muxOutConnector[38] = fifoOut[36][2];
              muxOutConnector[39] = fifoOut[37][2];
              muxOutConnector[40] = fifoOut[38][2];
              muxOutConnector[41] = fifoOut[39][2];
              muxOutConnector[42] = fifoOut[40][2];
              muxOutConnector[43] = fifoOut[41][2];
              muxOutConnector[44] = fifoOut[42][2];
              muxOutConnector[45] = fifoOut[43][2];
              muxOutConnector[46] = fifoOut[44][2];
              muxOutConnector[47] = fifoOut[45][2];
              muxOutConnector[48] = fifoOut[46][2];
              muxOutConnector[49] = fifoOut[47][2];
              muxOutConnector[50] = fifoOut[48][2];
              muxOutConnector[51] = fifoOut[49][2];
         end
         19: begin
              muxOutConnector[0] = fifoOut[19][9];
              muxOutConnector[1] = fifoOut[20][9];
              muxOutConnector[2] = fifoOut[21][9];
              muxOutConnector[3] = fifoOut[22][9];
              muxOutConnector[4] = fifoOut[23][9];
              muxOutConnector[5] = fifoOut[24][9];
              muxOutConnector[6] = fifoOut[25][9];
              muxOutConnector[7] = fifoOut[0][8];
              muxOutConnector[8] = fifoOut[1][8];
              muxOutConnector[9] = fifoOut[2][8];
              muxOutConnector[10] = fifoOut[3][8];
              muxOutConnector[11] = fifoOut[4][8];
              muxOutConnector[12] = fifoOut[5][8];
              muxOutConnector[13] = fifoOut[6][8];
              muxOutConnector[14] = fifoOut[7][8];
              muxOutConnector[15] = fifoOut[8][8];
              muxOutConnector[16] = fifoOut[9][8];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[50][2];
              muxOutConnector[27] = fifoOut[51][2];
              muxOutConnector[28] = fifoOut[26][1];
              muxOutConnector[29] = fifoOut[27][1];
              muxOutConnector[30] = fifoOut[28][1];
              muxOutConnector[31] = fifoOut[29][1];
              muxOutConnector[32] = fifoOut[30][1];
              muxOutConnector[33] = fifoOut[31][1];
              muxOutConnector[34] = fifoOut[32][1];
              muxOutConnector[35] = fifoOut[33][1];
              muxOutConnector[36] = fifoOut[34][1];
              muxOutConnector[37] = fifoOut[35][1];
              muxOutConnector[38] = fifoOut[36][1];
              muxOutConnector[39] = fifoOut[37][1];
              muxOutConnector[40] = fifoOut[38][1];
              muxOutConnector[41] = fifoOut[39][1];
              muxOutConnector[42] = fifoOut[40][1];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
         end
         default: begin
               for(i=0;i<muxOutSymbols;i=i+1)begin
                muxOutConnector[i] = 0;
              end
         end
//hgjhgbuiguigbigbgbgbui
         endcase
       case(rd_address_case)
         0: begin
              muxOutConnector_firstiter[0] = fifoOut[10][16];
              muxOutConnector_firstiter[1] = fifoOut[11][16];
              muxOutConnector_firstiter[2] = fifoOut[12][16];
              muxOutConnector_firstiter[3] = fifoOut[13][16];
              muxOutConnector_firstiter[4] = fifoOut[14][16];
              muxOutConnector_firstiter[5] = fifoOut[15][16];
              muxOutConnector_firstiter[6] = fifoOut[16][16];
              muxOutConnector_firstiter[7] = fifoOut[17][16];
              muxOutConnector_firstiter[8] = fifoOut[18][16];
              muxOutConnector_firstiter[9] = fifoOut[19][16];
              muxOutConnector_firstiter[10] = fifoOut[20][16];
              muxOutConnector_firstiter[11] = fifoOut[21][16];
              muxOutConnector_firstiter[12] = fifoOut[22][16];
              muxOutConnector_firstiter[13] = fifoOut[23][16];
              muxOutConnector_firstiter[14] = fifoOut[24][16];
              muxOutConnector_firstiter[15] = fifoOut[25][16];
              muxOutConnector_firstiter[16] = fifoOut[26][16];
              muxOutConnector_firstiter[17] = fifoOut[27][16];
              muxOutConnector_firstiter[18] = fifoOut[28][16];
              muxOutConnector_firstiter[19] = fifoOut[29][16];
              muxOutConnector_firstiter[20] = fifoOut[30][16];
              muxOutConnector_firstiter[21] = fifoOut[31][16];
              muxOutConnector_firstiter[22] = fifoOut[0][15];
              muxOutConnector_firstiter[23] = fifoOut[1][15];
              muxOutConnector_firstiter[24] = fifoOut[2][15];
              muxOutConnector_firstiter[25] = fifoOut[3][15];
              muxOutConnector_firstiter[26] = fifoOut[18][4];
              muxOutConnector_firstiter[27] = fifoOut[19][4];
              muxOutConnector_firstiter[28] = fifoOut[20][4];
              muxOutConnector_firstiter[29] = fifoOut[21][4];
              muxOutConnector_firstiter[30] = fifoOut[22][4];
              muxOutConnector_firstiter[31] = fifoOut[23][4];
              muxOutConnector_firstiter[32] = fifoOut[24][4];
              muxOutConnector_firstiter[33] = fifoOut[25][4];
              muxOutConnector_firstiter[34] = fifoOut[26][4];
              muxOutConnector_firstiter[35] = fifoOut[27][4];
              muxOutConnector_firstiter[36] = fifoOut[28][4];
              muxOutConnector_firstiter[37] = fifoOut[29][4];
              muxOutConnector_firstiter[38] = fifoOut[30][4];
              muxOutConnector_firstiter[39] = fifoOut[31][4];
              muxOutConnector_firstiter[40] = fifoOut[0][3];
              muxOutConnector_firstiter[41] = fifoOut[1][3];
              muxOutConnector_firstiter[42] = fifoOut[2][3];
              muxOutConnector_firstiter[43] = fifoOut[3][3];
              muxOutConnector_firstiter[44] = fifoOut[4][3];
              muxOutConnector_firstiter[45] = fifoOut[5][3];
              muxOutConnector_firstiter[46] = fifoOut[6][3];
              muxOutConnector_firstiter[47] = fifoOut[7][3];
              muxOutConnector_firstiter[48] = fifoOut[8][3];
              muxOutConnector_firstiter[49] = fifoOut[9][3];
              muxOutConnector_firstiter[50] = fifoOut[10][3];
              muxOutConnector_firstiter[51] = fifoOut[11][3];
         end
         1: begin
              muxOutConnector_firstiter[0] = fifoOut[4][15];
              muxOutConnector_firstiter[1] = fifoOut[5][15];
              muxOutConnector_firstiter[2] = fifoOut[6][15];
              muxOutConnector_firstiter[3] = fifoOut[7][15];
              muxOutConnector_firstiter[4] = fifoOut[8][15];
              muxOutConnector_firstiter[5] = fifoOut[9][15];
              muxOutConnector_firstiter[6] = fifoOut[10][15];
              muxOutConnector_firstiter[7] = fifoOut[11][15];
              muxOutConnector_firstiter[8] = fifoOut[12][15];
              muxOutConnector_firstiter[9] = fifoOut[13][15];
              muxOutConnector_firstiter[10] = fifoOut[14][15];
              muxOutConnector_firstiter[11] = fifoOut[15][15];
              muxOutConnector_firstiter[12] = fifoOut[16][15];
              muxOutConnector_firstiter[13] = fifoOut[17][15];
              muxOutConnector_firstiter[14] = fifoOut[18][15];
              muxOutConnector_firstiter[15] = fifoOut[19][15];
              muxOutConnector_firstiter[16] = fifoOut[20][15];
              muxOutConnector_firstiter[17] = fifoOut[21][15];
              muxOutConnector_firstiter[18] = fifoOut[22][15];
              muxOutConnector_firstiter[19] = fifoOut[23][15];
              muxOutConnector_firstiter[20] = fifoOut[24][15];
              muxOutConnector_firstiter[21] = fifoOut[25][15];
              muxOutConnector_firstiter[22] = fifoOut[26][15];
              muxOutConnector_firstiter[23] = fifoOut[27][15];
              muxOutConnector_firstiter[24] = fifoOut[28][15];
              muxOutConnector_firstiter[25] = fifoOut[29][15];
              muxOutConnector_firstiter[26] = fifoOut[12][3];
              muxOutConnector_firstiter[27] = fifoOut[13][3];
              muxOutConnector_firstiter[28] = fifoOut[14][3];
              muxOutConnector_firstiter[29] = fifoOut[15][3];
              muxOutConnector_firstiter[30] = fifoOut[16][3];
              muxOutConnector_firstiter[31] = fifoOut[17][3];
              muxOutConnector_firstiter[32] = fifoOut[18][3];
              muxOutConnector_firstiter[33] = fifoOut[19][3];
              muxOutConnector_firstiter[34] = fifoOut[20][3];
              muxOutConnector_firstiter[35] = fifoOut[21][3];
              muxOutConnector_firstiter[36] = fifoOut[22][3];
              muxOutConnector_firstiter[37] = fifoOut[23][3];
              muxOutConnector_firstiter[38] = fifoOut[24][3];
              muxOutConnector_firstiter[39] = fifoOut[25][3];
              muxOutConnector_firstiter[40] = fifoOut[26][3];
              muxOutConnector_firstiter[41] = fifoOut[27][3];
              muxOutConnector_firstiter[42] = fifoOut[28][3];
              muxOutConnector_firstiter[43] = fifoOut[29][3];
              muxOutConnector_firstiter[44] = fifoOut[30][3];
              muxOutConnector_firstiter[45] = fifoOut[31][3];
              muxOutConnector_firstiter[46] = fifoOut[0][2];
              muxOutConnector_firstiter[47] = fifoOut[1][2];
              muxOutConnector_firstiter[48] = fifoOut[2][2];
              muxOutConnector_firstiter[49] = fifoOut[3][2];
              muxOutConnector_firstiter[50] = fifoOut[4][2];
              muxOutConnector_firstiter[51] = fifoOut[5][2];
         end
         2: begin
              muxOutConnector_firstiter[0] = fifoOut[30][15];
              muxOutConnector_firstiter[1] = fifoOut[31][15];
              muxOutConnector_firstiter[2] = fifoOut[0][14];
              muxOutConnector_firstiter[3] = fifoOut[1][14];
              muxOutConnector_firstiter[4] = fifoOut[2][14];
              muxOutConnector_firstiter[5] = fifoOut[3][14];
              muxOutConnector_firstiter[6] = fifoOut[4][14];
              muxOutConnector_firstiter[7] = fifoOut[5][14];
              muxOutConnector_firstiter[8] = fifoOut[6][14];
              muxOutConnector_firstiter[9] = fifoOut[7][14];
              muxOutConnector_firstiter[10] = fifoOut[8][14];
              muxOutConnector_firstiter[11] = fifoOut[9][14];
              muxOutConnector_firstiter[12] = fifoOut[10][14];
              muxOutConnector_firstiter[13] = fifoOut[11][14];
              muxOutConnector_firstiter[14] = fifoOut[12][14];
              muxOutConnector_firstiter[15] = fifoOut[13][14];
              muxOutConnector_firstiter[16] = fifoOut[14][14];
              muxOutConnector_firstiter[17] = fifoOut[15][14];
              muxOutConnector_firstiter[18] = fifoOut[16][14];
              muxOutConnector_firstiter[19] = fifoOut[17][14];
              muxOutConnector_firstiter[20] = fifoOut[18][14];
              muxOutConnector_firstiter[21] = fifoOut[19][14];
              muxOutConnector_firstiter[22] = fifoOut[20][14];
              muxOutConnector_firstiter[23] = fifoOut[21][14];
              muxOutConnector_firstiter[24] = fifoOut[22][14];
              muxOutConnector_firstiter[25] = fifoOut[23][14];
              muxOutConnector_firstiter[26] = fifoOut[6][2];
              muxOutConnector_firstiter[27] = fifoOut[7][2];
              muxOutConnector_firstiter[28] = fifoOut[8][2];
              muxOutConnector_firstiter[29] = fifoOut[9][2];
              muxOutConnector_firstiter[30] = fifoOut[10][2];
              muxOutConnector_firstiter[31] = fifoOut[11][2];
              muxOutConnector_firstiter[32] = fifoOut[12][2];
              muxOutConnector_firstiter[33] = fifoOut[13][2];
              muxOutConnector_firstiter[34] = fifoOut[14][2];
              muxOutConnector_firstiter[35] = fifoOut[15][2];
              muxOutConnector_firstiter[36] = fifoOut[16][2];
              muxOutConnector_firstiter[37] = fifoOut[17][2];
              muxOutConnector_firstiter[38] = fifoOut[18][2];
              muxOutConnector_firstiter[39] = fifoOut[19][2];
              muxOutConnector_firstiter[40] = fifoOut[20][2];
              muxOutConnector_firstiter[41] = fifoOut[21][2];
              muxOutConnector_firstiter[42] = fifoOut[22][2];
              muxOutConnector_firstiter[43] = fifoOut[23][2];
              muxOutConnector_firstiter[44] = fifoOut[24][2];
              muxOutConnector_firstiter[45] = fifoOut[25][2];
              muxOutConnector_firstiter[46] = fifoOut[26][2];
              muxOutConnector_firstiter[47] = fifoOut[27][2];
              muxOutConnector_firstiter[48] = fifoOut[28][2];
              muxOutConnector_firstiter[49] = fifoOut[29][2];
              muxOutConnector_firstiter[50] = fifoOut[30][2];
              muxOutConnector_firstiter[51] = fifoOut[31][2];
         end
         3: begin
              muxOutConnector_firstiter[0] = fifoOut[24][14];
              muxOutConnector_firstiter[1] = fifoOut[25][14];
              muxOutConnector_firstiter[2] = fifoOut[26][14];
              muxOutConnector_firstiter[3] = fifoOut[27][14];
              muxOutConnector_firstiter[4] = fifoOut[28][14];
              muxOutConnector_firstiter[5] = fifoOut[29][14];
              muxOutConnector_firstiter[6] = fifoOut[30][14];
              muxOutConnector_firstiter[7] = fifoOut[31][14];
              muxOutConnector_firstiter[8] = fifoOut[0][13];
              muxOutConnector_firstiter[9] = fifoOut[1][13];
              muxOutConnector_firstiter[10] = fifoOut[2][13];
              muxOutConnector_firstiter[11] = fifoOut[3][13];
              muxOutConnector_firstiter[12] = fifoOut[4][13];
              muxOutConnector_firstiter[13] = fifoOut[5][13];
              muxOutConnector_firstiter[14] = fifoOut[6][13];
              muxOutConnector_firstiter[15] = fifoOut[7][13];
              muxOutConnector_firstiter[16] = fifoOut[8][13];
              muxOutConnector_firstiter[17] = fifoOut[9][13];
              muxOutConnector_firstiter[18] = fifoOut[10][13];
              muxOutConnector_firstiter[19] = fifoOut[11][13];
              muxOutConnector_firstiter[20] = fifoOut[12][13];
              muxOutConnector_firstiter[21] = fifoOut[13][13];
              muxOutConnector_firstiter[22] = fifoOut[14][13];
              muxOutConnector_firstiter[23] = fifoOut[15][13];
              muxOutConnector_firstiter[24] = fifoOut[16][13];
              muxOutConnector_firstiter[25] = fifoOut[17][13];
              muxOutConnector_firstiter[26] = fifoOut[0][1];
              muxOutConnector_firstiter[27] = fifoOut[1][1];
              muxOutConnector_firstiter[28] = fifoOut[2][1];
              muxOutConnector_firstiter[29] = fifoOut[3][1];
              muxOutConnector_firstiter[30] = fifoOut[4][1];
              muxOutConnector_firstiter[31] = fifoOut[5][1];
              muxOutConnector_firstiter[32] = fifoOut[6][1];
              muxOutConnector_firstiter[33] = fifoOut[7][1];
              muxOutConnector_firstiter[34] = fifoOut[8][1];
              muxOutConnector_firstiter[35] = fifoOut[9][1];
              muxOutConnector_firstiter[36] = fifoOut[10][1];
              muxOutConnector_firstiter[37] = fifoOut[11][1];
              muxOutConnector_firstiter[38] = fifoOut[12][1];
              muxOutConnector_firstiter[39] = fifoOut[13][1];
              muxOutConnector_firstiter[40] = fifoOut[14][1];
              muxOutConnector_firstiter[41] = fifoOut[15][1];
              muxOutConnector_firstiter[42] = fifoOut[16][1];
              muxOutConnector_firstiter[43] = fifoOut[17][1];
              muxOutConnector_firstiter[44] = fifoOut[18][1];
              muxOutConnector_firstiter[45] = fifoOut[19][1];
              muxOutConnector_firstiter[46] = fifoOut[20][1];
              muxOutConnector_firstiter[47] = fifoOut[21][1];
              muxOutConnector_firstiter[48] = fifoOut[22][1];
              muxOutConnector_firstiter[49] = fifoOut[23][1];
              muxOutConnector_firstiter[50] = fifoOut[24][1];
              muxOutConnector_firstiter[51] = fifoOut[25][1];
         end
         4: begin
              muxOutConnector_firstiter[0] = fifoOut[18][13];
              muxOutConnector_firstiter[1] = fifoOut[19][13];
              muxOutConnector_firstiter[2] = fifoOut[20][13];
              muxOutConnector_firstiter[3] = fifoOut[21][13];
              muxOutConnector_firstiter[4] = fifoOut[22][13];
              muxOutConnector_firstiter[5] = fifoOut[23][13];
              muxOutConnector_firstiter[6] = fifoOut[24][13];
              muxOutConnector_firstiter[7] = fifoOut[25][13];
              muxOutConnector_firstiter[8] = fifoOut[26][13];
              muxOutConnector_firstiter[9] = fifoOut[27][13];
              muxOutConnector_firstiter[10] = fifoOut[28][13];
              muxOutConnector_firstiter[11] = fifoOut[29][13];
              muxOutConnector_firstiter[12] = fifoOut[30][13];
              muxOutConnector_firstiter[13] = fifoOut[31][13];
              muxOutConnector_firstiter[14] = fifoOut[0][12];
              muxOutConnector_firstiter[15] = fifoOut[1][12];
              muxOutConnector_firstiter[16] = fifoOut[2][12];
              muxOutConnector_firstiter[17] = fifoOut[3][12];
              muxOutConnector_firstiter[18] = fifoOut[4][12];
              muxOutConnector_firstiter[19] = fifoOut[5][12];
              muxOutConnector_firstiter[20] = fifoOut[6][12];
              muxOutConnector_firstiter[21] = fifoOut[7][12];
              muxOutConnector_firstiter[22] = fifoOut[8][12];
              muxOutConnector_firstiter[23] = fifoOut[9][12];
              muxOutConnector_firstiter[24] = fifoOut[10][12];
              muxOutConnector_firstiter[25] = fifoOut[11][12];
              muxOutConnector_firstiter[26] = fifoOut[26][1];
              muxOutConnector_firstiter[27] = fifoOut[27][1];
              muxOutConnector_firstiter[28] = fifoOut[28][1];
              muxOutConnector_firstiter[29] = fifoOut[29][1];
              muxOutConnector_firstiter[30] = fifoOut[30][1];
              muxOutConnector_firstiter[31] = fifoOut[31][1];
              muxOutConnector_firstiter[32] = fifoOut[0][0];
              muxOutConnector_firstiter[33] = fifoOut[1][0];
              muxOutConnector_firstiter[34] = fifoOut[2][0];
              muxOutConnector_firstiter[35] = fifoOut[3][0];
              muxOutConnector_firstiter[36] = fifoOut[4][0];
              muxOutConnector_firstiter[37] = fifoOut[5][0];
              muxOutConnector_firstiter[38] = fifoOut[6][0];
              muxOutConnector_firstiter[39] = fifoOut[7][0];
              muxOutConnector_firstiter[40] = fifoOut[8][0];
              muxOutConnector_firstiter[41] = fifoOut[10][16];
              muxOutConnector_firstiter[42] = fifoOut[11][16];
              muxOutConnector_firstiter[43] = fifoOut[12][16];
              muxOutConnector_firstiter[44] = fifoOut[13][16];
              muxOutConnector_firstiter[45] = fifoOut[14][16];
              muxOutConnector_firstiter[46] = fifoOut[15][16];
              muxOutConnector_firstiter[47] = fifoOut[16][16];
              muxOutConnector_firstiter[48] = fifoOut[17][16];
              muxOutConnector_firstiter[49] = fifoOut[18][16];
              muxOutConnector_firstiter[50] = fifoOut[19][16];
              muxOutConnector_firstiter[51] = fifoOut[20][16];
         end
         5: begin
              muxOutConnector_firstiter[0] = fifoOut[12][12];
              muxOutConnector_firstiter[1] = fifoOut[13][12];
              muxOutConnector_firstiter[2] = fifoOut[14][12];
              muxOutConnector_firstiter[3] = fifoOut[15][12];
              muxOutConnector_firstiter[4] = fifoOut[16][12];
              muxOutConnector_firstiter[5] = fifoOut[17][12];
              muxOutConnector_firstiter[6] = fifoOut[18][12];
              muxOutConnector_firstiter[7] = fifoOut[19][12];
              muxOutConnector_firstiter[8] = fifoOut[20][12];
              muxOutConnector_firstiter[9] = fifoOut[21][12];
              muxOutConnector_firstiter[10] = fifoOut[22][12];
              muxOutConnector_firstiter[11] = fifoOut[23][12];
              muxOutConnector_firstiter[12] = fifoOut[24][12];
              muxOutConnector_firstiter[13] = fifoOut[25][12];
              muxOutConnector_firstiter[14] = fifoOut[26][12];
              muxOutConnector_firstiter[15] = fifoOut[27][12];
              muxOutConnector_firstiter[16] = fifoOut[28][12];
              muxOutConnector_firstiter[17] = fifoOut[29][12];
              muxOutConnector_firstiter[18] = fifoOut[30][12];
              muxOutConnector_firstiter[19] = fifoOut[31][12];
              muxOutConnector_firstiter[20] = fifoOut[0][11];
              muxOutConnector_firstiter[21] = fifoOut[1][11];
              muxOutConnector_firstiter[22] = fifoOut[2][11];
              muxOutConnector_firstiter[23] = fifoOut[3][11];
              muxOutConnector_firstiter[24] = fifoOut[4][11];
              muxOutConnector_firstiter[25] = fifoOut[5][11];
              muxOutConnector_firstiter[26] = fifoOut[21][16];
              muxOutConnector_firstiter[27] = fifoOut[22][16];
              muxOutConnector_firstiter[28] = fifoOut[23][16];
              muxOutConnector_firstiter[29] = fifoOut[24][16];
              muxOutConnector_firstiter[30] = fifoOut[25][16];
              muxOutConnector_firstiter[31] = fifoOut[26][16];
              muxOutConnector_firstiter[32] = fifoOut[27][16];
              muxOutConnector_firstiter[33] = fifoOut[28][16];
              muxOutConnector_firstiter[34] = fifoOut[29][16];
              muxOutConnector_firstiter[35] = fifoOut[30][16];
              muxOutConnector_firstiter[36] = fifoOut[31][16];
              muxOutConnector_firstiter[37] = fifoOut[0][15];
              muxOutConnector_firstiter[38] = fifoOut[1][15];
              muxOutConnector_firstiter[39] = fifoOut[2][15];
              muxOutConnector_firstiter[40] = fifoOut[3][15];
              muxOutConnector_firstiter[41] = fifoOut[4][15];
              muxOutConnector_firstiter[42] = fifoOut[5][15];
              muxOutConnector_firstiter[43] = fifoOut[6][15];
              muxOutConnector_firstiter[44] = fifoOut[7][15];
              muxOutConnector_firstiter[45] = fifoOut[8][15];
              muxOutConnector_firstiter[46] = fifoOut[9][15];
              muxOutConnector_firstiter[47] = fifoOut[10][15];
              muxOutConnector_firstiter[48] = fifoOut[11][15];
              muxOutConnector_firstiter[49] = fifoOut[12][15];
              muxOutConnector_firstiter[50] = fifoOut[13][15];
              muxOutConnector_firstiter[51] = fifoOut[14][15];
         end
         6: begin
              muxOutConnector_firstiter[0] = fifoOut[6][11];
              muxOutConnector_firstiter[1] = fifoOut[7][11];
              muxOutConnector_firstiter[2] = fifoOut[8][11];
              muxOutConnector_firstiter[3] = fifoOut[9][11];
              muxOutConnector_firstiter[4] = fifoOut[10][11];
              muxOutConnector_firstiter[5] = fifoOut[11][11];
              muxOutConnector_firstiter[6] = fifoOut[12][11];
              muxOutConnector_firstiter[7] = fifoOut[13][11];
              muxOutConnector_firstiter[8] = fifoOut[14][11];
              muxOutConnector_firstiter[9] = fifoOut[15][11];
              muxOutConnector_firstiter[10] = fifoOut[16][11];
              muxOutConnector_firstiter[11] = fifoOut[17][11];
              muxOutConnector_firstiter[12] = fifoOut[18][11];
              muxOutConnector_firstiter[13] = fifoOut[19][11];
              muxOutConnector_firstiter[14] = fifoOut[20][11];
              muxOutConnector_firstiter[15] = fifoOut[21][11];
              muxOutConnector_firstiter[16] = fifoOut[22][11];
              muxOutConnector_firstiter[17] = fifoOut[23][11];
              muxOutConnector_firstiter[18] = fifoOut[24][11];
              muxOutConnector_firstiter[19] = fifoOut[25][11];
              muxOutConnector_firstiter[20] = fifoOut[26][11];
              muxOutConnector_firstiter[21] = fifoOut[27][11];
              muxOutConnector_firstiter[22] = fifoOut[28][11];
              muxOutConnector_firstiter[23] = fifoOut[29][11];
              muxOutConnector_firstiter[24] = fifoOut[30][11];
              muxOutConnector_firstiter[25] = fifoOut[31][11];
              muxOutConnector_firstiter[26] = fifoOut[15][15];
              muxOutConnector_firstiter[27] = fifoOut[16][15];
              muxOutConnector_firstiter[28] = fifoOut[17][15];
              muxOutConnector_firstiter[29] = fifoOut[18][15];
              muxOutConnector_firstiter[30] = fifoOut[19][15];
              muxOutConnector_firstiter[31] = fifoOut[20][15];
              muxOutConnector_firstiter[32] = fifoOut[21][15];
              muxOutConnector_firstiter[33] = fifoOut[22][15];
              muxOutConnector_firstiter[34] = fifoOut[23][15];
              muxOutConnector_firstiter[35] = fifoOut[24][15];
              muxOutConnector_firstiter[36] = fifoOut[25][15];
              muxOutConnector_firstiter[37] = fifoOut[26][15];
              muxOutConnector_firstiter[38] = fifoOut[27][15];
              muxOutConnector_firstiter[39] = fifoOut[28][15];
              muxOutConnector_firstiter[40] = fifoOut[29][15];
              muxOutConnector_firstiter[41] = fifoOut[30][15];
              muxOutConnector_firstiter[42] = fifoOut[31][15];
              muxOutConnector_firstiter[43] = fifoOut[0][14];
              muxOutConnector_firstiter[44] = fifoOut[1][14];
              muxOutConnector_firstiter[45] = fifoOut[2][14];
              muxOutConnector_firstiter[46] = fifoOut[3][14];
              muxOutConnector_firstiter[47] = fifoOut[4][14];
              muxOutConnector_firstiter[48] = fifoOut[5][14];
              muxOutConnector_firstiter[49] = fifoOut[6][14];
              muxOutConnector_firstiter[50] = fifoOut[7][14];
              muxOutConnector_firstiter[51] = fifoOut[8][14];
         end
         7: begin
              muxOutConnector_firstiter[0] = fifoOut[0][10];
              muxOutConnector_firstiter[1] = fifoOut[1][10];
              muxOutConnector_firstiter[2] = fifoOut[2][10];
              muxOutConnector_firstiter[3] = fifoOut[3][10];
              muxOutConnector_firstiter[4] = fifoOut[4][10];
              muxOutConnector_firstiter[5] = fifoOut[5][10];
              muxOutConnector_firstiter[6] = fifoOut[6][10];
              muxOutConnector_firstiter[7] = fifoOut[7][10];
              muxOutConnector_firstiter[8] = fifoOut[8][10];
              muxOutConnector_firstiter[9] = fifoOut[9][10];
              muxOutConnector_firstiter[10] = fifoOut[10][10];
              muxOutConnector_firstiter[11] = fifoOut[11][10];
              muxOutConnector_firstiter[12] = fifoOut[12][10];
              muxOutConnector_firstiter[13] = fifoOut[13][10];
              muxOutConnector_firstiter[14] = fifoOut[14][10];
              muxOutConnector_firstiter[15] = fifoOut[15][10];
              muxOutConnector_firstiter[16] = fifoOut[16][10];
              muxOutConnector_firstiter[17] = fifoOut[17][10];
              muxOutConnector_firstiter[18] = fifoOut[18][10];
              muxOutConnector_firstiter[19] = fifoOut[19][10];
              muxOutConnector_firstiter[20] = fifoOut[20][10];
              muxOutConnector_firstiter[21] = fifoOut[21][10];
              muxOutConnector_firstiter[22] = fifoOut[22][10];
              muxOutConnector_firstiter[23] = fifoOut[23][10];
              muxOutConnector_firstiter[24] = fifoOut[24][10];
              muxOutConnector_firstiter[25] = fifoOut[25][10];
              muxOutConnector_firstiter[26] = fifoOut[9][14];
              muxOutConnector_firstiter[27] = fifoOut[10][14];
              muxOutConnector_firstiter[28] = fifoOut[11][14];
              muxOutConnector_firstiter[29] = fifoOut[12][14];
              muxOutConnector_firstiter[30] = fifoOut[13][14];
              muxOutConnector_firstiter[31] = fifoOut[14][14];
              muxOutConnector_firstiter[32] = fifoOut[15][14];
              muxOutConnector_firstiter[33] = fifoOut[16][14];
              muxOutConnector_firstiter[34] = fifoOut[17][14];
              muxOutConnector_firstiter[35] = fifoOut[18][14];
              muxOutConnector_firstiter[36] = fifoOut[19][14];
              muxOutConnector_firstiter[37] = fifoOut[20][14];
              muxOutConnector_firstiter[38] = fifoOut[21][14];
              muxOutConnector_firstiter[39] = fifoOut[22][14];
              muxOutConnector_firstiter[40] = fifoOut[23][14];
              muxOutConnector_firstiter[41] = fifoOut[24][14];
              muxOutConnector_firstiter[42] = fifoOut[25][14];
              muxOutConnector_firstiter[43] = fifoOut[26][14];
              muxOutConnector_firstiter[44] = fifoOut[27][14];
              muxOutConnector_firstiter[45] = fifoOut[28][14];
              muxOutConnector_firstiter[46] = fifoOut[29][14];
              muxOutConnector_firstiter[47] = fifoOut[30][14];
              muxOutConnector_firstiter[48] = fifoOut[31][14];
              muxOutConnector_firstiter[49] = fifoOut[0][13];
              muxOutConnector_firstiter[50] = fifoOut[1][13];
              muxOutConnector_firstiter[51] = fifoOut[2][13];
         end
         8: begin
              muxOutConnector_firstiter[0] = fifoOut[26][10];
              muxOutConnector_firstiter[1] = fifoOut[27][10];
              muxOutConnector_firstiter[2] = fifoOut[28][10];
              muxOutConnector_firstiter[3] = fifoOut[29][10];
              muxOutConnector_firstiter[4] = fifoOut[30][10];
              muxOutConnector_firstiter[5] = fifoOut[31][10];
              muxOutConnector_firstiter[6] = fifoOut[0][9];
              muxOutConnector_firstiter[7] = fifoOut[1][9];
              muxOutConnector_firstiter[8] = fifoOut[2][9];
              muxOutConnector_firstiter[9] = fifoOut[3][9];
              muxOutConnector_firstiter[10] = fifoOut[4][9];
              muxOutConnector_firstiter[11] = fifoOut[5][9];
              muxOutConnector_firstiter[12] = fifoOut[6][9];
              muxOutConnector_firstiter[13] = fifoOut[7][9];
              muxOutConnector_firstiter[14] = fifoOut[8][9];
              muxOutConnector_firstiter[15] = fifoOut[9][9];
              muxOutConnector_firstiter[16] = fifoOut[10][9];
              muxOutConnector_firstiter[17] = fifoOut[11][9];
              muxOutConnector_firstiter[18] = fifoOut[12][9];
              muxOutConnector_firstiter[19] = fifoOut[13][9];
              muxOutConnector_firstiter[20] = fifoOut[14][9];
              muxOutConnector_firstiter[21] = fifoOut[15][9];
              muxOutConnector_firstiter[22] = fifoOut[16][9];
              muxOutConnector_firstiter[23] = fifoOut[17][9];
              muxOutConnector_firstiter[24] = fifoOut[18][9];
              muxOutConnector_firstiter[25] = fifoOut[19][9];
              muxOutConnector_firstiter[26] = fifoOut[3][13];
              muxOutConnector_firstiter[27] = fifoOut[4][13];
              muxOutConnector_firstiter[28] = fifoOut[5][13];
              muxOutConnector_firstiter[29] = fifoOut[6][13];
              muxOutConnector_firstiter[30] = fifoOut[7][13];
              muxOutConnector_firstiter[31] = fifoOut[8][13];
              muxOutConnector_firstiter[32] = fifoOut[9][13];
              muxOutConnector_firstiter[33] = fifoOut[10][13];
              muxOutConnector_firstiter[34] = fifoOut[11][13];
              muxOutConnector_firstiter[35] = fifoOut[12][13];
              muxOutConnector_firstiter[36] = fifoOut[13][13];
              muxOutConnector_firstiter[37] = fifoOut[14][13];
              muxOutConnector_firstiter[38] = fifoOut[15][13];
              muxOutConnector_firstiter[39] = fifoOut[16][13];
              muxOutConnector_firstiter[40] = fifoOut[17][13];
              muxOutConnector_firstiter[41] = fifoOut[18][13];
              muxOutConnector_firstiter[42] = fifoOut[19][13];
              muxOutConnector_firstiter[43] = fifoOut[20][13];
              muxOutConnector_firstiter[44] = fifoOut[21][13];
              muxOutConnector_firstiter[45] = fifoOut[22][13];
              muxOutConnector_firstiter[46] = fifoOut[23][13];
              muxOutConnector_firstiter[47] = fifoOut[24][13];
              muxOutConnector_firstiter[48] = fifoOut[25][13];
              muxOutConnector_firstiter[49] = fifoOut[26][13];
              muxOutConnector_firstiter[50] = fifoOut[27][13];
              muxOutConnector_firstiter[51] = fifoOut[28][13];
         end
         9: begin
              muxOutConnector_firstiter[0] = fifoOut[20][9];
              muxOutConnector_firstiter[1] = fifoOut[21][9];
              muxOutConnector_firstiter[2] = fifoOut[22][9];
              muxOutConnector_firstiter[3] = fifoOut[23][9];
              muxOutConnector_firstiter[4] = fifoOut[24][9];
              muxOutConnector_firstiter[5] = fifoOut[25][9];
              muxOutConnector_firstiter[6] = fifoOut[26][9];
              muxOutConnector_firstiter[7] = fifoOut[27][9];
              muxOutConnector_firstiter[8] = fifoOut[28][9];
              muxOutConnector_firstiter[9] = fifoOut[29][9];
              muxOutConnector_firstiter[10] = fifoOut[30][9];
              muxOutConnector_firstiter[11] = fifoOut[31][9];
              muxOutConnector_firstiter[12] = fifoOut[0][8];
              muxOutConnector_firstiter[13] = fifoOut[1][8];
              muxOutConnector_firstiter[14] = fifoOut[2][8];
              muxOutConnector_firstiter[15] = fifoOut[3][8];
              muxOutConnector_firstiter[16] = fifoOut[4][8];
              muxOutConnector_firstiter[17] = fifoOut[5][8];
              muxOutConnector_firstiter[18] = fifoOut[6][8];
              muxOutConnector_firstiter[19] = fifoOut[7][8];
              muxOutConnector_firstiter[20] = fifoOut[8][8];
              muxOutConnector_firstiter[21] = fifoOut[9][8];
              muxOutConnector_firstiter[22] = fifoOut[10][8];
              muxOutConnector_firstiter[23] = fifoOut[11][8];
              muxOutConnector_firstiter[24] = fifoOut[12][8];
              muxOutConnector_firstiter[25] = fifoOut[13][8];
              muxOutConnector_firstiter[26] = fifoOut[29][13];
              muxOutConnector_firstiter[27] = fifoOut[30][13];
              muxOutConnector_firstiter[28] = fifoOut[31][13];
              muxOutConnector_firstiter[29] = fifoOut[0][12];
              muxOutConnector_firstiter[30] = fifoOut[1][12];
              muxOutConnector_firstiter[31] = fifoOut[2][12];
              muxOutConnector_firstiter[32] = fifoOut[3][12];
              muxOutConnector_firstiter[33] = fifoOut[4][12];
              muxOutConnector_firstiter[34] = fifoOut[5][12];
              muxOutConnector_firstiter[35] = fifoOut[6][12];
              muxOutConnector_firstiter[36] = fifoOut[7][12];
              muxOutConnector_firstiter[37] = fifoOut[8][12];
              muxOutConnector_firstiter[38] = fifoOut[9][12];
              muxOutConnector_firstiter[39] = fifoOut[10][12];
              muxOutConnector_firstiter[40] = fifoOut[11][12];
              muxOutConnector_firstiter[41] = fifoOut[12][12];
              muxOutConnector_firstiter[42] = fifoOut[13][12];
              muxOutConnector_firstiter[43] = fifoOut[14][12];
              muxOutConnector_firstiter[44] = fifoOut[15][12];
              muxOutConnector_firstiter[45] = fifoOut[16][12];
              muxOutConnector_firstiter[46] = fifoOut[17][12];
              muxOutConnector_firstiter[47] = fifoOut[18][12];
              muxOutConnector_firstiter[48] = fifoOut[19][12];
              muxOutConnector_firstiter[49] = fifoOut[20][12];
              muxOutConnector_firstiter[50] = fifoOut[21][12];
              muxOutConnector_firstiter[51] = fifoOut[22][12];
         end
         10: begin
              muxOutConnector_firstiter[0] = fifoOut[14][8];
              muxOutConnector_firstiter[1] = fifoOut[15][8];
              muxOutConnector_firstiter[2] = fifoOut[16][8];
              muxOutConnector_firstiter[3] = fifoOut[17][8];
              muxOutConnector_firstiter[4] = fifoOut[18][8];
              muxOutConnector_firstiter[5] = fifoOut[19][8];
              muxOutConnector_firstiter[6] = fifoOut[20][8];
              muxOutConnector_firstiter[7] = fifoOut[21][8];
              muxOutConnector_firstiter[8] = fifoOut[22][8];
              muxOutConnector_firstiter[9] = fifoOut[23][8];
              muxOutConnector_firstiter[10] = fifoOut[24][8];
              muxOutConnector_firstiter[11] = fifoOut[25][8];
              muxOutConnector_firstiter[12] = fifoOut[26][8];
              muxOutConnector_firstiter[13] = fifoOut[27][8];
              muxOutConnector_firstiter[14] = fifoOut[28][8];
              muxOutConnector_firstiter[15] = fifoOut[29][8];
              muxOutConnector_firstiter[16] = fifoOut[30][8];
              muxOutConnector_firstiter[17] = fifoOut[31][8];
              muxOutConnector_firstiter[18] = fifoOut[0][7];
              muxOutConnector_firstiter[19] = fifoOut[1][7];
              muxOutConnector_firstiter[20] = fifoOut[2][7];
              muxOutConnector_firstiter[21] = fifoOut[3][7];
              muxOutConnector_firstiter[22] = fifoOut[4][7];
              muxOutConnector_firstiter[23] = fifoOut[5][7];
              muxOutConnector_firstiter[24] = fifoOut[6][7];
              muxOutConnector_firstiter[25] = fifoOut[7][7];
              muxOutConnector_firstiter[26] = fifoOut[23][12];
              muxOutConnector_firstiter[27] = fifoOut[24][12];
              muxOutConnector_firstiter[28] = fifoOut[25][12];
              muxOutConnector_firstiter[29] = fifoOut[26][12];
              muxOutConnector_firstiter[30] = fifoOut[27][12];
              muxOutConnector_firstiter[31] = fifoOut[28][12];
              muxOutConnector_firstiter[32] = fifoOut[29][12];
              muxOutConnector_firstiter[33] = fifoOut[30][12];
              muxOutConnector_firstiter[34] = fifoOut[31][12];
              muxOutConnector_firstiter[35] = fifoOut[0][11];
              muxOutConnector_firstiter[36] = fifoOut[1][11];
              muxOutConnector_firstiter[37] = fifoOut[2][11];
              muxOutConnector_firstiter[38] = fifoOut[3][11];
              muxOutConnector_firstiter[39] = fifoOut[4][11];
              muxOutConnector_firstiter[40] = fifoOut[5][11];
              muxOutConnector_firstiter[41] = fifoOut[6][11];
              muxOutConnector_firstiter[42] = fifoOut[7][11];
              muxOutConnector_firstiter[43] = fifoOut[8][11];
              muxOutConnector_firstiter[44] = fifoOut[9][11];
              muxOutConnector_firstiter[45] = fifoOut[10][11];
              muxOutConnector_firstiter[46] = fifoOut[11][11];
              muxOutConnector_firstiter[47] = fifoOut[12][11];
              muxOutConnector_firstiter[48] = fifoOut[13][11];
              muxOutConnector_firstiter[49] = fifoOut[14][11];
              muxOutConnector_firstiter[50] = fifoOut[15][11];
              muxOutConnector_firstiter[51] = fifoOut[16][11];
         end
         11: begin
              muxOutConnector_firstiter[0] = fifoOut[8][7];
              muxOutConnector_firstiter[1] = fifoOut[9][7];
              muxOutConnector_firstiter[2] = fifoOut[10][7];
              muxOutConnector_firstiter[3] = fifoOut[11][7];
              muxOutConnector_firstiter[4] = fifoOut[12][7];
              muxOutConnector_firstiter[5] = fifoOut[13][7];
              muxOutConnector_firstiter[6] = fifoOut[14][7];
              muxOutConnector_firstiter[7] = fifoOut[15][7];
              muxOutConnector_firstiter[8] = fifoOut[16][7];
              muxOutConnector_firstiter[9] = fifoOut[17][7];
              muxOutConnector_firstiter[10] = fifoOut[18][7];
              muxOutConnector_firstiter[11] = fifoOut[19][7];
              muxOutConnector_firstiter[12] = fifoOut[20][7];
              muxOutConnector_firstiter[13] = fifoOut[21][7];
              muxOutConnector_firstiter[14] = fifoOut[22][7];
              muxOutConnector_firstiter[15] = fifoOut[23][7];
              muxOutConnector_firstiter[16] = fifoOut[24][7];
              muxOutConnector_firstiter[17] = fifoOut[25][7];
              muxOutConnector_firstiter[18] = fifoOut[26][7];
              muxOutConnector_firstiter[19] = fifoOut[27][7];
              muxOutConnector_firstiter[20] = fifoOut[28][7];
              muxOutConnector_firstiter[21] = fifoOut[29][7];
              muxOutConnector_firstiter[22] = fifoOut[30][7];
              muxOutConnector_firstiter[23] = fifoOut[31][7];
              muxOutConnector_firstiter[24] = fifoOut[0][6];
              muxOutConnector_firstiter[25] = fifoOut[1][6];
              muxOutConnector_firstiter[26] = fifoOut[17][11];
              muxOutConnector_firstiter[27] = fifoOut[18][11];
              muxOutConnector_firstiter[28] = fifoOut[19][11];
              muxOutConnector_firstiter[29] = fifoOut[20][11];
              muxOutConnector_firstiter[30] = fifoOut[21][11];
              muxOutConnector_firstiter[31] = fifoOut[22][11];
              muxOutConnector_firstiter[32] = fifoOut[23][11];
              muxOutConnector_firstiter[33] = fifoOut[24][11];
              muxOutConnector_firstiter[34] = fifoOut[25][11];
              muxOutConnector_firstiter[35] = fifoOut[26][11];
              muxOutConnector_firstiter[36] = fifoOut[27][11];
              muxOutConnector_firstiter[37] = fifoOut[28][11];
              muxOutConnector_firstiter[38] = fifoOut[29][11];
              muxOutConnector_firstiter[39] = fifoOut[30][11];
              muxOutConnector_firstiter[40] = fifoOut[31][11];
              muxOutConnector_firstiter[41] = fifoOut[0][10];
              muxOutConnector_firstiter[42] = fifoOut[1][10];
              muxOutConnector_firstiter[43] = fifoOut[2][10];
              muxOutConnector_firstiter[44] = fifoOut[3][10];
              muxOutConnector_firstiter[45] = fifoOut[4][10];
              muxOutConnector_firstiter[46] = fifoOut[5][10];
              muxOutConnector_firstiter[47] = fifoOut[6][10];
              muxOutConnector_firstiter[48] = fifoOut[7][10];
              muxOutConnector_firstiter[49] = fifoOut[8][10];
              muxOutConnector_firstiter[50] = fifoOut[9][10];
              muxOutConnector_firstiter[51] = fifoOut[10][10];
         end
         12: begin
              muxOutConnector_firstiter[0] = fifoOut[2][6];
              muxOutConnector_firstiter[1] = fifoOut[3][6];
              muxOutConnector_firstiter[2] = fifoOut[4][6];
              muxOutConnector_firstiter[3] = fifoOut[5][6];
              muxOutConnector_firstiter[4] = fifoOut[6][6];
              muxOutConnector_firstiter[5] = fifoOut[7][6];
              muxOutConnector_firstiter[6] = fifoOut[8][6];
              muxOutConnector_firstiter[7] = fifoOut[9][6];
              muxOutConnector_firstiter[8] = fifoOut[10][6];
              muxOutConnector_firstiter[9] = fifoOut[11][6];
              muxOutConnector_firstiter[10] = fifoOut[12][6];
              muxOutConnector_firstiter[11] = fifoOut[13][6];
              muxOutConnector_firstiter[12] = fifoOut[14][6];
              muxOutConnector_firstiter[13] = fifoOut[15][6];
              muxOutConnector_firstiter[14] = fifoOut[16][6];
              muxOutConnector_firstiter[15] = fifoOut[17][6];
              muxOutConnector_firstiter[16] = fifoOut[18][6];
              muxOutConnector_firstiter[17] = fifoOut[19][6];
              muxOutConnector_firstiter[18] = fifoOut[20][6];
              muxOutConnector_firstiter[19] = fifoOut[21][6];
              muxOutConnector_firstiter[20] = fifoOut[22][6];
              muxOutConnector_firstiter[21] = fifoOut[23][6];
              muxOutConnector_firstiter[22] = fifoOut[24][6];
              muxOutConnector_firstiter[23] = fifoOut[25][6];
              muxOutConnector_firstiter[24] = fifoOut[26][6];
              muxOutConnector_firstiter[25] = fifoOut[27][6];
              muxOutConnector_firstiter[26] = fifoOut[11][10];
              muxOutConnector_firstiter[27] = fifoOut[12][10];
              muxOutConnector_firstiter[28] = fifoOut[13][10];
              muxOutConnector_firstiter[29] = fifoOut[14][10];
              muxOutConnector_firstiter[30] = fifoOut[15][10];
              muxOutConnector_firstiter[31] = fifoOut[16][10];
              muxOutConnector_firstiter[32] = fifoOut[17][10];
              muxOutConnector_firstiter[33] = fifoOut[18][10];
              muxOutConnector_firstiter[34] = fifoOut[19][10];
              muxOutConnector_firstiter[35] = fifoOut[20][10];
              muxOutConnector_firstiter[36] = fifoOut[21][10];
              muxOutConnector_firstiter[37] = fifoOut[22][10];
              muxOutConnector_firstiter[38] = fifoOut[23][10];
              muxOutConnector_firstiter[39] = fifoOut[24][10];
              muxOutConnector_firstiter[40] = fifoOut[25][10];
              muxOutConnector_firstiter[41] = fifoOut[26][10];
              muxOutConnector_firstiter[42] = fifoOut[27][10];
              muxOutConnector_firstiter[43] = fifoOut[28][10];
              muxOutConnector_firstiter[44] = fifoOut[29][10];
              muxOutConnector_firstiter[45] = fifoOut[30][10];
              muxOutConnector_firstiter[46] = fifoOut[31][10];
              muxOutConnector_firstiter[47] = fifoOut[0][9];
              muxOutConnector_firstiter[48] = fifoOut[1][9];
              muxOutConnector_firstiter[49] = fifoOut[2][9];
              muxOutConnector_firstiter[50] = fifoOut[3][9];
              muxOutConnector_firstiter[51] = fifoOut[4][9];
         end
         13: begin
              muxOutConnector_firstiter[0] = fifoOut[28][6];
              muxOutConnector_firstiter[1] = fifoOut[29][6];
              muxOutConnector_firstiter[2] = fifoOut[30][6];
              muxOutConnector_firstiter[3] = fifoOut[31][6];
              muxOutConnector_firstiter[4] = fifoOut[0][5];
              muxOutConnector_firstiter[5] = fifoOut[1][5];
              muxOutConnector_firstiter[6] = fifoOut[2][5];
              muxOutConnector_firstiter[7] = fifoOut[3][5];
              muxOutConnector_firstiter[8] = fifoOut[4][5];
              muxOutConnector_firstiter[9] = fifoOut[5][5];
              muxOutConnector_firstiter[10] = fifoOut[6][5];
              muxOutConnector_firstiter[11] = fifoOut[7][5];
              muxOutConnector_firstiter[12] = fifoOut[8][5];
              muxOutConnector_firstiter[13] = fifoOut[9][5];
              muxOutConnector_firstiter[14] = fifoOut[10][5];
              muxOutConnector_firstiter[15] = fifoOut[11][5];
              muxOutConnector_firstiter[16] = fifoOut[12][5];
              muxOutConnector_firstiter[17] = fifoOut[13][5];
              muxOutConnector_firstiter[18] = fifoOut[14][5];
              muxOutConnector_firstiter[19] = fifoOut[15][5];
              muxOutConnector_firstiter[20] = fifoOut[16][5];
              muxOutConnector_firstiter[21] = fifoOut[17][5];
              muxOutConnector_firstiter[22] = fifoOut[18][5];
              muxOutConnector_firstiter[23] = fifoOut[19][5];
              muxOutConnector_firstiter[24] = fifoOut[20][5];
              muxOutConnector_firstiter[25] = fifoOut[21][5];
              muxOutConnector_firstiter[26] = fifoOut[5][9];
              muxOutConnector_firstiter[27] = fifoOut[6][9];
              muxOutConnector_firstiter[28] = fifoOut[7][9];
              muxOutConnector_firstiter[29] = fifoOut[8][9];
              muxOutConnector_firstiter[30] = fifoOut[9][9];
              muxOutConnector_firstiter[31] = fifoOut[10][9];
              muxOutConnector_firstiter[32] = fifoOut[11][9];
              muxOutConnector_firstiter[33] = fifoOut[12][9];
              muxOutConnector_firstiter[34] = fifoOut[13][9];
              muxOutConnector_firstiter[35] = fifoOut[14][9];
              muxOutConnector_firstiter[36] = fifoOut[15][9];
              muxOutConnector_firstiter[37] = fifoOut[16][9];
              muxOutConnector_firstiter[38] = fifoOut[17][9];
              muxOutConnector_firstiter[39] = fifoOut[18][9];
              muxOutConnector_firstiter[40] = fifoOut[19][9];
              muxOutConnector_firstiter[41] = fifoOut[20][9];
              muxOutConnector_firstiter[42] = fifoOut[21][9];
              muxOutConnector_firstiter[43] = fifoOut[22][9];
              muxOutConnector_firstiter[44] = fifoOut[23][9];
              muxOutConnector_firstiter[45] = fifoOut[24][9];
              muxOutConnector_firstiter[46] = fifoOut[25][9];
              muxOutConnector_firstiter[47] = fifoOut[26][9];
              muxOutConnector_firstiter[48] = fifoOut[27][9];
              muxOutConnector_firstiter[49] = fifoOut[28][9];
              muxOutConnector_firstiter[50] = fifoOut[29][9];
              muxOutConnector_firstiter[51] = fifoOut[30][9];
         end
         14: begin
              muxOutConnector_firstiter[0] = fifoOut[22][5];
              muxOutConnector_firstiter[1] = fifoOut[23][5];
              muxOutConnector_firstiter[2] = fifoOut[24][5];
              muxOutConnector_firstiter[3] = fifoOut[25][5];
              muxOutConnector_firstiter[4] = fifoOut[26][5];
              muxOutConnector_firstiter[5] = fifoOut[27][5];
              muxOutConnector_firstiter[6] = fifoOut[28][5];
              muxOutConnector_firstiter[7] = fifoOut[29][5];
              muxOutConnector_firstiter[8] = fifoOut[30][5];
              muxOutConnector_firstiter[9] = fifoOut[31][5];
              muxOutConnector_firstiter[10] = fifoOut[0][4];
              muxOutConnector_firstiter[11] = fifoOut[1][4];
              muxOutConnector_firstiter[12] = fifoOut[2][4];
              muxOutConnector_firstiter[13] = fifoOut[3][4];
              muxOutConnector_firstiter[14] = fifoOut[4][4];
              muxOutConnector_firstiter[15] = fifoOut[5][4];
              muxOutConnector_firstiter[16] = fifoOut[6][4];
              muxOutConnector_firstiter[17] = fifoOut[7][4];
              muxOutConnector_firstiter[18] = fifoOut[8][4];
              muxOutConnector_firstiter[19] = fifoOut[9][4];
              muxOutConnector_firstiter[20] = fifoOut[10][4];
              muxOutConnector_firstiter[21] = fifoOut[11][4];
              muxOutConnector_firstiter[22] = fifoOut[12][4];
              muxOutConnector_firstiter[23] = fifoOut[13][4];
              muxOutConnector_firstiter[24] = fifoOut[14][4];
              muxOutConnector_firstiter[25] = fifoOut[15][4];
              muxOutConnector_firstiter[26] = fifoOut[31][9];
              muxOutConnector_firstiter[27] = fifoOut[0][8];
              muxOutConnector_firstiter[28] = fifoOut[1][8];
              muxOutConnector_firstiter[29] = fifoOut[2][8];
              muxOutConnector_firstiter[30] = fifoOut[3][8];
              muxOutConnector_firstiter[31] = fifoOut[4][8];
              muxOutConnector_firstiter[32] = fifoOut[5][8];
              muxOutConnector_firstiter[33] = fifoOut[6][8];
              muxOutConnector_firstiter[34] = fifoOut[7][8];
              muxOutConnector_firstiter[35] = fifoOut[8][8];
              muxOutConnector_firstiter[36] = fifoOut[9][8];
              muxOutConnector_firstiter[37] = fifoOut[10][8];
              muxOutConnector_firstiter[38] = fifoOut[11][8];
              muxOutConnector_firstiter[39] = fifoOut[12][8];
              muxOutConnector_firstiter[40] = fifoOut[13][8];
              muxOutConnector_firstiter[41] = fifoOut[14][8];
              muxOutConnector_firstiter[42] = fifoOut[15][8];
              muxOutConnector_firstiter[43] = fifoOut[16][8];
              muxOutConnector_firstiter[44] = fifoOut[17][8];
              muxOutConnector_firstiter[45] = fifoOut[18][8];
              muxOutConnector_firstiter[46] = fifoOut[19][8];
              muxOutConnector_firstiter[47] = fifoOut[20][8];
              muxOutConnector_firstiter[48] = fifoOut[21][8];
              muxOutConnector_firstiter[49] = fifoOut[22][8];
              muxOutConnector_firstiter[50] = fifoOut[23][8];
              muxOutConnector_firstiter[51] = fifoOut[24][8];
         end
         15: begin
              muxOutConnector_firstiter[0] = fifoOut[16][4];
              muxOutConnector_firstiter[1] = fifoOut[17][4];
              muxOutConnector_firstiter[2] = fifoOut[18][4];
              muxOutConnector_firstiter[3] = fifoOut[19][4];
              muxOutConnector_firstiter[4] = fifoOut[20][4];
              muxOutConnector_firstiter[5] = fifoOut[21][4];
              muxOutConnector_firstiter[6] = fifoOut[22][4];
              muxOutConnector_firstiter[7] = fifoOut[23][4];
              muxOutConnector_firstiter[8] = fifoOut[24][4];
              muxOutConnector_firstiter[9] = fifoOut[25][4];
              muxOutConnector_firstiter[10] = fifoOut[26][4];
              muxOutConnector_firstiter[11] = fifoOut[27][4];
              muxOutConnector_firstiter[12] = fifoOut[28][4];
              muxOutConnector_firstiter[13] = fifoOut[29][4];
              muxOutConnector_firstiter[14] = fifoOut[30][4];
              muxOutConnector_firstiter[15] = fifoOut[31][4];
              muxOutConnector_firstiter[16] = fifoOut[0][3];
              muxOutConnector_firstiter[17] = fifoOut[1][3];
              muxOutConnector_firstiter[18] = fifoOut[2][3];
              muxOutConnector_firstiter[19] = fifoOut[3][3];
              muxOutConnector_firstiter[20] = fifoOut[4][3];
              muxOutConnector_firstiter[21] = fifoOut[5][3];
              muxOutConnector_firstiter[22] = fifoOut[6][3];
              muxOutConnector_firstiter[23] = fifoOut[7][3];
              muxOutConnector_firstiter[24] = fifoOut[8][3];
              muxOutConnector_firstiter[25] = fifoOut[9][3];
              muxOutConnector_firstiter[26] = fifoOut[25][8];
              muxOutConnector_firstiter[27] = fifoOut[26][8];
              muxOutConnector_firstiter[28] = fifoOut[27][8];
              muxOutConnector_firstiter[29] = fifoOut[28][8];
              muxOutConnector_firstiter[30] = fifoOut[29][8];
              muxOutConnector_firstiter[31] = fifoOut[30][8];
              muxOutConnector_firstiter[32] = fifoOut[31][8];
              muxOutConnector_firstiter[33] = fifoOut[0][7];
              muxOutConnector_firstiter[34] = fifoOut[1][7];
              muxOutConnector_firstiter[35] = fifoOut[2][7];
              muxOutConnector_firstiter[36] = fifoOut[3][7];
              muxOutConnector_firstiter[37] = fifoOut[4][7];
              muxOutConnector_firstiter[38] = fifoOut[5][7];
              muxOutConnector_firstiter[39] = fifoOut[6][7];
              muxOutConnector_firstiter[40] = fifoOut[7][7];
              muxOutConnector_firstiter[41] = fifoOut[8][7];
              muxOutConnector_firstiter[42] = fifoOut[9][7];
              muxOutConnector_firstiter[43] = fifoOut[10][7];
              muxOutConnector_firstiter[44] = fifoOut[11][7];
              muxOutConnector_firstiter[45] = fifoOut[12][7];
              muxOutConnector_firstiter[46] = fifoOut[13][7];
              muxOutConnector_firstiter[47] = fifoOut[14][7];
              muxOutConnector_firstiter[48] = fifoOut[15][7];
              muxOutConnector_firstiter[49] = fifoOut[16][7];
              muxOutConnector_firstiter[50] = fifoOut[17][7];
              muxOutConnector_firstiter[51] = fifoOut[18][7];
         end
         16: begin
              muxOutConnector_firstiter[0] = fifoOut[10][3];
              muxOutConnector_firstiter[1] = fifoOut[11][3];
              muxOutConnector_firstiter[2] = fifoOut[12][3];
              muxOutConnector_firstiter[3] = fifoOut[13][3];
              muxOutConnector_firstiter[4] = fifoOut[14][3];
              muxOutConnector_firstiter[5] = fifoOut[15][3];
              muxOutConnector_firstiter[6] = fifoOut[16][3];
              muxOutConnector_firstiter[7] = fifoOut[17][3];
              muxOutConnector_firstiter[8] = fifoOut[18][3];
              muxOutConnector_firstiter[9] = fifoOut[19][3];
              muxOutConnector_firstiter[10] = fifoOut[20][3];
              muxOutConnector_firstiter[11] = fifoOut[21][3];
              muxOutConnector_firstiter[12] = fifoOut[22][3];
              muxOutConnector_firstiter[13] = fifoOut[23][3];
              muxOutConnector_firstiter[14] = fifoOut[24][3];
              muxOutConnector_firstiter[15] = fifoOut[25][3];
              muxOutConnector_firstiter[16] = fifoOut[26][3];
              muxOutConnector_firstiter[17] = fifoOut[27][3];
              muxOutConnector_firstiter[18] = fifoOut[28][3];
              muxOutConnector_firstiter[19] = fifoOut[29][3];
              muxOutConnector_firstiter[20] = fifoOut[30][3];
              muxOutConnector_firstiter[21] = fifoOut[31][3];
              muxOutConnector_firstiter[22] = fifoOut[0][2];
              muxOutConnector_firstiter[23] = fifoOut[1][2];
              muxOutConnector_firstiter[24] = fifoOut[2][2];
              muxOutConnector_firstiter[25] = fifoOut[3][2];
              muxOutConnector_firstiter[26] = fifoOut[19][7];
              muxOutConnector_firstiter[27] = fifoOut[20][7];
              muxOutConnector_firstiter[28] = fifoOut[21][7];
              muxOutConnector_firstiter[29] = fifoOut[22][7];
              muxOutConnector_firstiter[30] = fifoOut[23][7];
              muxOutConnector_firstiter[31] = fifoOut[24][7];
              muxOutConnector_firstiter[32] = fifoOut[25][7];
              muxOutConnector_firstiter[33] = fifoOut[26][7];
              muxOutConnector_firstiter[34] = fifoOut[27][7];
              muxOutConnector_firstiter[35] = fifoOut[28][7];
              muxOutConnector_firstiter[36] = fifoOut[29][7];
              muxOutConnector_firstiter[37] = fifoOut[30][7];
              muxOutConnector_firstiter[38] = fifoOut[31][7];
              muxOutConnector_firstiter[39] = fifoOut[0][6];
              muxOutConnector_firstiter[40] = fifoOut[1][6];
              muxOutConnector_firstiter[41] = fifoOut[2][6];
              muxOutConnector_firstiter[42] = fifoOut[3][6];
              muxOutConnector_firstiter[43] = fifoOut[4][6];
              muxOutConnector_firstiter[44] = fifoOut[5][6];
              muxOutConnector_firstiter[45] = fifoOut[6][6];
              muxOutConnector_firstiter[46] = fifoOut[7][6];
              muxOutConnector_firstiter[47] = fifoOut[8][6];
              muxOutConnector_firstiter[48] = fifoOut[9][6];
              muxOutConnector_firstiter[49] = fifoOut[10][6];
              muxOutConnector_firstiter[50] = fifoOut[11][6];
              muxOutConnector_firstiter[51] = fifoOut[12][6];
         end
         17: begin
              muxOutConnector_firstiter[0] = fifoOut[4][2];
              muxOutConnector_firstiter[1] = fifoOut[5][2];
              muxOutConnector_firstiter[2] = fifoOut[6][2];
              muxOutConnector_firstiter[3] = fifoOut[7][2];
              muxOutConnector_firstiter[4] = fifoOut[8][2];
              muxOutConnector_firstiter[5] = fifoOut[9][2];
              muxOutConnector_firstiter[6] = fifoOut[10][2];
              muxOutConnector_firstiter[7] = fifoOut[11][2];
              muxOutConnector_firstiter[8] = fifoOut[12][2];
              muxOutConnector_firstiter[9] = fifoOut[13][2];
              muxOutConnector_firstiter[10] = fifoOut[14][2];
              muxOutConnector_firstiter[11] = fifoOut[15][2];
              muxOutConnector_firstiter[12] = fifoOut[16][2];
              muxOutConnector_firstiter[13] = fifoOut[17][2];
              muxOutConnector_firstiter[14] = fifoOut[18][2];
              muxOutConnector_firstiter[15] = fifoOut[19][2];
              muxOutConnector_firstiter[16] = fifoOut[20][2];
              muxOutConnector_firstiter[17] = fifoOut[21][2];
              muxOutConnector_firstiter[18] = fifoOut[22][2];
              muxOutConnector_firstiter[19] = fifoOut[23][2];
              muxOutConnector_firstiter[20] = fifoOut[24][2];
              muxOutConnector_firstiter[21] = fifoOut[25][2];
              muxOutConnector_firstiter[22] = fifoOut[26][2];
              muxOutConnector_firstiter[23] = fifoOut[27][2];
              muxOutConnector_firstiter[24] = fifoOut[28][2];
              muxOutConnector_firstiter[25] = fifoOut[29][2];
              muxOutConnector_firstiter[26] = fifoOut[13][6];
              muxOutConnector_firstiter[27] = fifoOut[14][6];
              muxOutConnector_firstiter[28] = fifoOut[15][6];
              muxOutConnector_firstiter[29] = fifoOut[16][6];
              muxOutConnector_firstiter[30] = fifoOut[17][6];
              muxOutConnector_firstiter[31] = fifoOut[18][6];
              muxOutConnector_firstiter[32] = fifoOut[19][6];
              muxOutConnector_firstiter[33] = fifoOut[20][6];
              muxOutConnector_firstiter[34] = fifoOut[21][6];
              muxOutConnector_firstiter[35] = fifoOut[22][6];
              muxOutConnector_firstiter[36] = fifoOut[23][6];
              muxOutConnector_firstiter[37] = fifoOut[24][6];
              muxOutConnector_firstiter[38] = fifoOut[25][6];
              muxOutConnector_firstiter[39] = fifoOut[26][6];
              muxOutConnector_firstiter[40] = fifoOut[27][6];
              muxOutConnector_firstiter[41] = fifoOut[28][6];
              muxOutConnector_firstiter[42] = fifoOut[29][6];
              muxOutConnector_firstiter[43] = fifoOut[30][6];
              muxOutConnector_firstiter[44] = fifoOut[31][6];
              muxOutConnector_firstiter[45] = fifoOut[0][5];
              muxOutConnector_firstiter[46] = fifoOut[1][5];
              muxOutConnector_firstiter[47] = fifoOut[2][5];
              muxOutConnector_firstiter[48] = fifoOut[3][5];
              muxOutConnector_firstiter[49] = fifoOut[4][5];
              muxOutConnector_firstiter[50] = fifoOut[5][5];
              muxOutConnector_firstiter[51] = fifoOut[6][5];
         end
         18: begin
              muxOutConnector_firstiter[0] = fifoOut[30][2];
              muxOutConnector_firstiter[1] = fifoOut[31][2];
              muxOutConnector_firstiter[2] = fifoOut[0][1];
              muxOutConnector_firstiter[3] = fifoOut[1][1];
              muxOutConnector_firstiter[4] = fifoOut[2][1];
              muxOutConnector_firstiter[5] = fifoOut[3][1];
              muxOutConnector_firstiter[6] = fifoOut[4][1];
              muxOutConnector_firstiter[7] = fifoOut[5][1];
              muxOutConnector_firstiter[8] = fifoOut[6][1];
              muxOutConnector_firstiter[9] = fifoOut[7][1];
              muxOutConnector_firstiter[10] = fifoOut[8][1];
              muxOutConnector_firstiter[11] = fifoOut[9][1];
              muxOutConnector_firstiter[12] = fifoOut[10][1];
              muxOutConnector_firstiter[13] = fifoOut[11][1];
              muxOutConnector_firstiter[14] = fifoOut[12][1];
              muxOutConnector_firstiter[15] = fifoOut[13][1];
              muxOutConnector_firstiter[16] = fifoOut[14][1];
              muxOutConnector_firstiter[17] = fifoOut[15][1];
              muxOutConnector_firstiter[18] = fifoOut[16][1];
              muxOutConnector_firstiter[19] = fifoOut[17][1];
              muxOutConnector_firstiter[20] = fifoOut[18][1];
              muxOutConnector_firstiter[21] = fifoOut[19][1];
              muxOutConnector_firstiter[22] = fifoOut[20][1];
              muxOutConnector_firstiter[23] = fifoOut[21][1];
              muxOutConnector_firstiter[24] = fifoOut[22][1];
              muxOutConnector_firstiter[25] = fifoOut[23][1];
              muxOutConnector_firstiter[26] = fifoOut[7][5];
              muxOutConnector_firstiter[27] = fifoOut[8][5];
              muxOutConnector_firstiter[28] = fifoOut[9][5];
              muxOutConnector_firstiter[29] = fifoOut[10][5];
              muxOutConnector_firstiter[30] = fifoOut[11][5];
              muxOutConnector_firstiter[31] = fifoOut[12][5];
              muxOutConnector_firstiter[32] = fifoOut[13][5];
              muxOutConnector_firstiter[33] = fifoOut[14][5];
              muxOutConnector_firstiter[34] = fifoOut[15][5];
              muxOutConnector_firstiter[35] = fifoOut[16][5];
              muxOutConnector_firstiter[36] = fifoOut[17][5];
              muxOutConnector_firstiter[37] = fifoOut[18][5];
              muxOutConnector_firstiter[38] = fifoOut[19][5];
              muxOutConnector_firstiter[39] = fifoOut[20][5];
              muxOutConnector_firstiter[40] = fifoOut[21][5];
              muxOutConnector_firstiter[41] = fifoOut[22][5];
              muxOutConnector_firstiter[42] = fifoOut[23][5];
              muxOutConnector_firstiter[43] = fifoOut[24][5];
              muxOutConnector_firstiter[44] = fifoOut[25][5];
              muxOutConnector_firstiter[45] = fifoOut[26][5];
              muxOutConnector_firstiter[46] = fifoOut[27][5];
              muxOutConnector_firstiter[47] = fifoOut[28][5];
              muxOutConnector_firstiter[48] = fifoOut[29][5];
              muxOutConnector_firstiter[49] = fifoOut[30][5];
              muxOutConnector_firstiter[50] = fifoOut[31][5];
              muxOutConnector_firstiter[51] = fifoOut[0][4];
         end
         19: begin
              muxOutConnector_firstiter[0] = fifoOut[24][1];
              muxOutConnector_firstiter[1] = fifoOut[25][1];
              muxOutConnector_firstiter[2] = fifoOut[26][1];
              muxOutConnector_firstiter[3] = fifoOut[27][1];
              muxOutConnector_firstiter[4] = fifoOut[28][1];
              muxOutConnector_firstiter[5] = fifoOut[29][1];
              muxOutConnector_firstiter[6] = fifoOut[30][1];
              muxOutConnector_firstiter[7] = fifoOut[31][1];
              muxOutConnector_firstiter[8] = fifoOut[0][0];
              muxOutConnector_firstiter[9] = fifoOut[1][0];
              muxOutConnector_firstiter[10] = fifoOut[2][0];
              muxOutConnector_firstiter[11] = fifoOut[3][0];
              muxOutConnector_firstiter[12] = fifoOut[4][0];
              muxOutConnector_firstiter[13] = fifoOut[5][0];
              muxOutConnector_firstiter[14] = fifoOut[6][0];
              muxOutConnector_firstiter[15] = fifoOut[7][0];
              muxOutConnector_firstiter[16] = fifoOut[8][0];
              muxOutConnector_firstiter[17] = maxVal;
              muxOutConnector_firstiter[18] = maxVal;
              muxOutConnector_firstiter[19] = maxVal;
              muxOutConnector_firstiter[20] = maxVal;
              muxOutConnector_firstiter[21] = maxVal;
              muxOutConnector_firstiter[22] = maxVal;
              muxOutConnector_firstiter[23] = maxVal;
              muxOutConnector_firstiter[24] = maxVal;
              muxOutConnector_firstiter[25] = maxVal;
              muxOutConnector_firstiter[26] = fifoOut[1][4];
              muxOutConnector_firstiter[27] = fifoOut[2][4];
              muxOutConnector_firstiter[28] = fifoOut[3][4];
              muxOutConnector_firstiter[29] = fifoOut[4][4];
              muxOutConnector_firstiter[30] = fifoOut[5][4];
              muxOutConnector_firstiter[31] = fifoOut[6][4];
              muxOutConnector_firstiter[32] = fifoOut[7][4];
              muxOutConnector_firstiter[33] = fifoOut[8][4];
              muxOutConnector_firstiter[34] = fifoOut[9][4];
              muxOutConnector_firstiter[35] = fifoOut[10][4];
              muxOutConnector_firstiter[36] = fifoOut[11][4];
              muxOutConnector_firstiter[37] = fifoOut[12][4];
              muxOutConnector_firstiter[38] = fifoOut[13][4];
              muxOutConnector_firstiter[39] = fifoOut[14][4];
              muxOutConnector_firstiter[40] = fifoOut[15][4];
              muxOutConnector_firstiter[41] = fifoOut[16][4];
              muxOutConnector_firstiter[42] = fifoOut[17][4];
              muxOutConnector_firstiter[43] = maxVal;
              muxOutConnector_firstiter[44] = maxVal;
              muxOutConnector_firstiter[45] = maxVal;
              muxOutConnector_firstiter[46] = maxVal;
              muxOutConnector_firstiter[47] = maxVal;
              muxOutConnector_firstiter[48] = maxVal;
              muxOutConnector_firstiter[49] = maxVal;
              muxOutConnector_firstiter[50] = maxVal;
              muxOutConnector_firstiter[51] = maxVal;
         end
         default: begin
               for(i=0;i<muxOutSymbols;i=i+1)begin
                muxOutConnector_firstiter[i] = 0;
              end
         end
     endcase
end//always
endmodule
