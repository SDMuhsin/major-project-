`timescale 1ns / 1ps
module LMem0To1_511_circ3_ys_scripted(
        muxOut,
        ly0In,
        wr_en,
        feedback_en,
        rd_address,
        rd_en,
        clk,
        rst
);
input feedback_en;
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 16;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        if(feedback_en) begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= fifoOut[i][c-1];
         end
        end
        else begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= ly0InConnector[i];
         end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[2][10];
              muxOutConnector[1] = fifoOut[3][10];
              muxOutConnector[2] = fifoOut[4][10];
              muxOutConnector[3] = fifoOut[5][10];
              muxOutConnector[4] = fifoOut[6][10];
              muxOutConnector[5] = fifoOut[7][10];
              muxOutConnector[6] = fifoOut[8][10];
              muxOutConnector[7] = fifoOut[9][10];
              muxOutConnector[8] = fifoOut[10][10];
              muxOutConnector[9] = fifoOut[11][10];
              muxOutConnector[10] = fifoOut[12][10];
              muxOutConnector[11] = fifoOut[13][10];
              muxOutConnector[12] = fifoOut[14][10];
              muxOutConnector[13] = fifoOut[15][10];
              muxOutConnector[14] = fifoOut[16][10];
              muxOutConnector[15] = fifoOut[17][10];
              muxOutConnector[16] = fifoOut[18][10];
              muxOutConnector[17] = fifoOut[19][10];
              muxOutConnector[18] = fifoOut[20][10];
              muxOutConnector[19] = fifoOut[21][10];
              muxOutConnector[20] = fifoOut[22][10];
              muxOutConnector[21] = fifoOut[23][10];
              muxOutConnector[22] = fifoOut[24][10];
              muxOutConnector[23] = fifoOut[25][10];
              muxOutConnector[24] = fifoOut[0][9];
              muxOutConnector[25] = fifoOut[1][9];
              muxOutConnector[26] = fifoOut[12][2];
              muxOutConnector[27] = fifoOut[13][2];
              muxOutConnector[28] = fifoOut[14][2];
              muxOutConnector[29] = fifoOut[15][2];
              muxOutConnector[30] = fifoOut[16][2];
              muxOutConnector[31] = fifoOut[17][2];
              muxOutConnector[32] = fifoOut[18][2];
              muxOutConnector[33] = fifoOut[19][2];
              muxOutConnector[34] = fifoOut[20][2];
              muxOutConnector[35] = fifoOut[21][2];
              muxOutConnector[36] = fifoOut[22][2];
              muxOutConnector[37] = fifoOut[23][2];
              muxOutConnector[38] = fifoOut[24][2];
              muxOutConnector[39] = fifoOut[25][2];
              muxOutConnector[40] = fifoOut[0][1];
              muxOutConnector[41] = fifoOut[1][1];
              muxOutConnector[42] = fifoOut[2][1];
              muxOutConnector[43] = fifoOut[3][1];
              muxOutConnector[44] = fifoOut[4][1];
              muxOutConnector[45] = fifoOut[5][1];
              muxOutConnector[46] = fifoOut[6][1];
              muxOutConnector[47] = fifoOut[7][1];
              muxOutConnector[48] = fifoOut[8][1];
              muxOutConnector[49] = fifoOut[9][1];
              muxOutConnector[50] = fifoOut[10][1];
              muxOutConnector[51] = fifoOut[11][1];
       end
       1: begin
              muxOutConnector[0] = fifoOut[2][10];
              muxOutConnector[1] = fifoOut[3][10];
              muxOutConnector[2] = fifoOut[4][10];
              muxOutConnector[3] = fifoOut[5][10];
              muxOutConnector[4] = fifoOut[6][10];
              muxOutConnector[5] = fifoOut[7][10];
              muxOutConnector[6] = fifoOut[8][10];
              muxOutConnector[7] = fifoOut[9][10];
              muxOutConnector[8] = fifoOut[10][10];
              muxOutConnector[9] = fifoOut[11][10];
              muxOutConnector[10] = fifoOut[12][10];
              muxOutConnector[11] = fifoOut[13][10];
              muxOutConnector[12] = fifoOut[14][10];
              muxOutConnector[13] = fifoOut[15][10];
              muxOutConnector[14] = fifoOut[16][10];
              muxOutConnector[15] = fifoOut[17][10];
              muxOutConnector[16] = fifoOut[18][10];
              muxOutConnector[17] = fifoOut[19][10];
              muxOutConnector[18] = fifoOut[20][10];
              muxOutConnector[19] = fifoOut[21][10];
              muxOutConnector[20] = fifoOut[22][10];
              muxOutConnector[21] = fifoOut[23][10];
              muxOutConnector[22] = fifoOut[24][10];
              muxOutConnector[23] = fifoOut[25][10];
              muxOutConnector[24] = fifoOut[0][9];
              muxOutConnector[25] = fifoOut[1][9];
              muxOutConnector[26] = fifoOut[12][2];
              muxOutConnector[27] = fifoOut[13][2];
              muxOutConnector[28] = fifoOut[14][2];
              muxOutConnector[29] = fifoOut[15][2];
              muxOutConnector[30] = fifoOut[16][2];
              muxOutConnector[31] = fifoOut[17][2];
              muxOutConnector[32] = fifoOut[18][2];
              muxOutConnector[33] = fifoOut[19][2];
              muxOutConnector[34] = fifoOut[20][2];
              muxOutConnector[35] = fifoOut[21][2];
              muxOutConnector[36] = fifoOut[22][2];
              muxOutConnector[37] = fifoOut[23][2];
              muxOutConnector[38] = fifoOut[24][2];
              muxOutConnector[39] = fifoOut[25][2];
              muxOutConnector[40] = fifoOut[0][1];
              muxOutConnector[41] = fifoOut[1][1];
              muxOutConnector[42] = fifoOut[2][1];
              muxOutConnector[43] = fifoOut[3][1];
              muxOutConnector[44] = fifoOut[4][1];
              muxOutConnector[45] = fifoOut[5][1];
              muxOutConnector[46] = fifoOut[6][1];
              muxOutConnector[47] = fifoOut[7][1];
              muxOutConnector[48] = fifoOut[8][1];
              muxOutConnector[49] = fifoOut[9][1];
              muxOutConnector[50] = fifoOut[10][1];
              muxOutConnector[51] = fifoOut[11][1];
       end
       2: begin
              muxOutConnector[0] = fifoOut[2][10];
              muxOutConnector[1] = fifoOut[3][10];
              muxOutConnector[2] = fifoOut[4][10];
              muxOutConnector[3] = fifoOut[5][10];
              muxOutConnector[4] = fifoOut[6][10];
              muxOutConnector[5] = fifoOut[7][10];
              muxOutConnector[6] = fifoOut[8][10];
              muxOutConnector[7] = fifoOut[9][10];
              muxOutConnector[8] = fifoOut[10][10];
              muxOutConnector[9] = fifoOut[11][10];
              muxOutConnector[10] = fifoOut[12][10];
              muxOutConnector[11] = fifoOut[13][10];
              muxOutConnector[12] = fifoOut[14][10];
              muxOutConnector[13] = fifoOut[15][10];
              muxOutConnector[14] = fifoOut[16][10];
              muxOutConnector[15] = fifoOut[17][10];
              muxOutConnector[16] = fifoOut[18][10];
              muxOutConnector[17] = fifoOut[19][10];
              muxOutConnector[18] = fifoOut[20][10];
              muxOutConnector[19] = fifoOut[21][10];
              muxOutConnector[20] = fifoOut[22][10];
              muxOutConnector[21] = fifoOut[23][10];
              muxOutConnector[22] = fifoOut[24][10];
              muxOutConnector[23] = fifoOut[25][10];
              muxOutConnector[24] = fifoOut[0][9];
              muxOutConnector[25] = fifoOut[1][9];
              muxOutConnector[26] = fifoOut[12][2];
              muxOutConnector[27] = fifoOut[13][2];
              muxOutConnector[28] = fifoOut[14][2];
              muxOutConnector[29] = fifoOut[15][2];
              muxOutConnector[30] = fifoOut[16][2];
              muxOutConnector[31] = fifoOut[26][1];
              muxOutConnector[32] = fifoOut[27][1];
              muxOutConnector[33] = fifoOut[28][1];
              muxOutConnector[34] = fifoOut[29][1];
              muxOutConnector[35] = fifoOut[30][1];
              muxOutConnector[36] = fifoOut[31][1];
              muxOutConnector[37] = fifoOut[32][1];
              muxOutConnector[38] = fifoOut[33][1];
              muxOutConnector[39] = fifoOut[34][1];
              muxOutConnector[40] = fifoOut[35][1];
              muxOutConnector[41] = fifoOut[36][1];
              muxOutConnector[42] = fifoOut[37][1];
              muxOutConnector[43] = fifoOut[38][1];
              muxOutConnector[44] = fifoOut[39][1];
              muxOutConnector[45] = fifoOut[40][1];
              muxOutConnector[46] = fifoOut[41][1];
              muxOutConnector[47] = fifoOut[42][1];
              muxOutConnector[48] = fifoOut[43][1];
              muxOutConnector[49] = fifoOut[44][1];
              muxOutConnector[50] = fifoOut[45][1];
              muxOutConnector[51] = fifoOut[46][1];
       end
       3: begin
              muxOutConnector[0] = fifoOut[2][10];
              muxOutConnector[1] = fifoOut[3][10];
              muxOutConnector[2] = fifoOut[4][10];
              muxOutConnector[3] = fifoOut[5][10];
              muxOutConnector[4] = fifoOut[6][10];
              muxOutConnector[5] = fifoOut[7][10];
              muxOutConnector[6] = fifoOut[8][10];
              muxOutConnector[7] = fifoOut[9][10];
              muxOutConnector[8] = fifoOut[10][10];
              muxOutConnector[9] = fifoOut[11][10];
              muxOutConnector[10] = fifoOut[12][10];
              muxOutConnector[11] = fifoOut[13][10];
              muxOutConnector[12] = fifoOut[14][10];
              muxOutConnector[13] = fifoOut[15][10];
              muxOutConnector[14] = fifoOut[16][10];
              muxOutConnector[15] = fifoOut[17][10];
              muxOutConnector[16] = fifoOut[18][10];
              muxOutConnector[17] = fifoOut[19][10];
              muxOutConnector[18] = fifoOut[20][10];
              muxOutConnector[19] = fifoOut[21][10];
              muxOutConnector[20] = fifoOut[22][10];
              muxOutConnector[21] = fifoOut[23][10];
              muxOutConnector[22] = fifoOut[24][10];
              muxOutConnector[23] = fifoOut[25][10];
              muxOutConnector[24] = fifoOut[0][9];
              muxOutConnector[25] = fifoOut[1][9];
              muxOutConnector[26] = fifoOut[47][2];
              muxOutConnector[27] = fifoOut[48][2];
              muxOutConnector[28] = fifoOut[49][2];
              muxOutConnector[29] = fifoOut[50][2];
              muxOutConnector[30] = fifoOut[51][2];
              muxOutConnector[31] = fifoOut[26][1];
              muxOutConnector[32] = fifoOut[27][1];
              muxOutConnector[33] = fifoOut[28][1];
              muxOutConnector[34] = fifoOut[29][1];
              muxOutConnector[35] = fifoOut[30][1];
              muxOutConnector[36] = fifoOut[31][1];
              muxOutConnector[37] = fifoOut[32][1];
              muxOutConnector[38] = fifoOut[33][1];
              muxOutConnector[39] = fifoOut[34][1];
              muxOutConnector[40] = fifoOut[35][1];
              muxOutConnector[41] = fifoOut[36][1];
              muxOutConnector[42] = fifoOut[37][1];
              muxOutConnector[43] = fifoOut[38][1];
              muxOutConnector[44] = fifoOut[39][1];
              muxOutConnector[45] = fifoOut[40][1];
              muxOutConnector[46] = fifoOut[41][1];
              muxOutConnector[47] = fifoOut[42][1];
              muxOutConnector[48] = fifoOut[43][1];
              muxOutConnector[49] = fifoOut[44][1];
              muxOutConnector[50] = fifoOut[45][1];
              muxOutConnector[51] = fifoOut[46][1];
       end
       4: begin
              muxOutConnector[0] = fifoOut[2][10];
              muxOutConnector[1] = fifoOut[3][10];
              muxOutConnector[2] = fifoOut[4][10];
              muxOutConnector[3] = fifoOut[5][10];
              muxOutConnector[4] = fifoOut[6][10];
              muxOutConnector[5] = fifoOut[7][10];
              muxOutConnector[6] = fifoOut[8][10];
              muxOutConnector[7] = fifoOut[9][10];
              muxOutConnector[8] = fifoOut[10][10];
              muxOutConnector[9] = fifoOut[11][10];
              muxOutConnector[10] = fifoOut[12][10];
              muxOutConnector[11] = fifoOut[13][10];
              muxOutConnector[12] = fifoOut[14][10];
              muxOutConnector[13] = fifoOut[15][10];
              muxOutConnector[14] = fifoOut[16][10];
              muxOutConnector[15] = fifoOut[17][10];
              muxOutConnector[16] = fifoOut[18][10];
              muxOutConnector[17] = fifoOut[19][10];
              muxOutConnector[18] = fifoOut[20][10];
              muxOutConnector[19] = fifoOut[21][10];
              muxOutConnector[20] = fifoOut[22][10];
              muxOutConnector[21] = fifoOut[23][10];
              muxOutConnector[22] = fifoOut[24][10];
              muxOutConnector[23] = fifoOut[25][10];
              muxOutConnector[24] = fifoOut[0][9];
              muxOutConnector[25] = fifoOut[1][9];
              muxOutConnector[26] = fifoOut[47][2];
              muxOutConnector[27] = fifoOut[48][2];
              muxOutConnector[28] = fifoOut[49][2];
              muxOutConnector[29] = fifoOut[50][2];
              muxOutConnector[30] = fifoOut[51][2];
              muxOutConnector[31] = fifoOut[26][1];
              muxOutConnector[32] = fifoOut[27][1];
              muxOutConnector[33] = fifoOut[28][1];
              muxOutConnector[34] = fifoOut[29][1];
              muxOutConnector[35] = fifoOut[30][1];
              muxOutConnector[36] = fifoOut[31][1];
              muxOutConnector[37] = fifoOut[32][1];
              muxOutConnector[38] = fifoOut[33][1];
              muxOutConnector[39] = fifoOut[34][1];
              muxOutConnector[40] = fifoOut[35][1];
              muxOutConnector[41] = fifoOut[36][1];
              muxOutConnector[42] = fifoOut[37][1];
              muxOutConnector[43] = fifoOut[38][1];
              muxOutConnector[44] = fifoOut[39][1];
              muxOutConnector[45] = fifoOut[40][1];
              muxOutConnector[46] = fifoOut[41][1];
              muxOutConnector[47] = fifoOut[42][1];
              muxOutConnector[48] = fifoOut[43][1];
              muxOutConnector[49] = fifoOut[44][1];
              muxOutConnector[50] = fifoOut[45][1];
              muxOutConnector[51] = fifoOut[46][1];
       end
       5: begin
              muxOutConnector[0] = fifoOut[2][10];
              muxOutConnector[1] = fifoOut[3][10];
              muxOutConnector[2] = fifoOut[4][10];
              muxOutConnector[3] = fifoOut[5][10];
              muxOutConnector[4] = fifoOut[6][10];
              muxOutConnector[5] = fifoOut[7][10];
              muxOutConnector[6] = fifoOut[8][10];
              muxOutConnector[7] = fifoOut[9][10];
              muxOutConnector[8] = fifoOut[10][10];
              muxOutConnector[9] = fifoOut[11][10];
              muxOutConnector[10] = fifoOut[12][10];
              muxOutConnector[11] = fifoOut[13][10];
              muxOutConnector[12] = fifoOut[14][10];
              muxOutConnector[13] = fifoOut[15][10];
              muxOutConnector[14] = fifoOut[16][10];
              muxOutConnector[15] = fifoOut[17][10];
              muxOutConnector[16] = fifoOut[18][10];
              muxOutConnector[17] = fifoOut[19][10];
              muxOutConnector[18] = fifoOut[20][10];
              muxOutConnector[19] = fifoOut[21][10];
              muxOutConnector[20] = fifoOut[22][10];
              muxOutConnector[21] = fifoOut[23][10];
              muxOutConnector[22] = fifoOut[24][10];
              muxOutConnector[23] = fifoOut[25][10];
              muxOutConnector[24] = fifoOut[0][9];
              muxOutConnector[25] = fifoOut[1][9];
              muxOutConnector[26] = fifoOut[47][2];
              muxOutConnector[27] = fifoOut[48][2];
              muxOutConnector[28] = fifoOut[49][2];
              muxOutConnector[29] = fifoOut[50][2];
              muxOutConnector[30] = fifoOut[51][2];
              muxOutConnector[31] = fifoOut[26][1];
              muxOutConnector[32] = fifoOut[27][1];
              muxOutConnector[33] = fifoOut[28][1];
              muxOutConnector[34] = fifoOut[29][1];
              muxOutConnector[35] = fifoOut[30][1];
              muxOutConnector[36] = fifoOut[31][1];
              muxOutConnector[37] = fifoOut[32][1];
              muxOutConnector[38] = fifoOut[33][1];
              muxOutConnector[39] = fifoOut[34][1];
              muxOutConnector[40] = fifoOut[35][1];
              muxOutConnector[41] = fifoOut[36][1];
              muxOutConnector[42] = fifoOut[37][1];
              muxOutConnector[43] = fifoOut[38][1];
              muxOutConnector[44] = fifoOut[39][1];
              muxOutConnector[45] = fifoOut[40][1];
              muxOutConnector[46] = fifoOut[41][1];
              muxOutConnector[47] = fifoOut[42][1];
              muxOutConnector[48] = fifoOut[43][1];
              muxOutConnector[49] = fifoOut[44][1];
              muxOutConnector[50] = fifoOut[45][1];
              muxOutConnector[51] = fifoOut[46][1];
       end
       6: begin
              muxOutConnector[0] = fifoOut[2][10];
              muxOutConnector[1] = fifoOut[3][10];
              muxOutConnector[2] = fifoOut[4][10];
              muxOutConnector[3] = fifoOut[5][10];
              muxOutConnector[4] = fifoOut[6][10];
              muxOutConnector[5] = fifoOut[7][10];
              muxOutConnector[6] = fifoOut[8][10];
              muxOutConnector[7] = fifoOut[9][10];
              muxOutConnector[8] = fifoOut[10][10];
              muxOutConnector[9] = fifoOut[11][10];
              muxOutConnector[10] = fifoOut[12][10];
              muxOutConnector[11] = fifoOut[13][10];
              muxOutConnector[12] = fifoOut[14][10];
              muxOutConnector[13] = fifoOut[15][10];
              muxOutConnector[14] = fifoOut[16][10];
              muxOutConnector[15] = fifoOut[17][10];
              muxOutConnector[16] = fifoOut[18][10];
              muxOutConnector[17] = fifoOut[19][10];
              muxOutConnector[18] = fifoOut[20][10];
              muxOutConnector[19] = fifoOut[21][10];
              muxOutConnector[20] = fifoOut[22][10];
              muxOutConnector[21] = fifoOut[23][10];
              muxOutConnector[22] = fifoOut[24][10];
              muxOutConnector[23] = fifoOut[25][10];
              muxOutConnector[24] = fifoOut[0][9];
              muxOutConnector[25] = fifoOut[1][9];
              muxOutConnector[26] = fifoOut[47][2];
              muxOutConnector[27] = fifoOut[48][2];
              muxOutConnector[28] = fifoOut[49][2];
              muxOutConnector[29] = fifoOut[50][2];
              muxOutConnector[30] = fifoOut[51][2];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = fifoOut[12][5];
              muxOutConnector[44] = fifoOut[13][5];
              muxOutConnector[45] = fifoOut[14][5];
              muxOutConnector[46] = fifoOut[15][5];
              muxOutConnector[47] = fifoOut[16][5];
              muxOutConnector[48] = fifoOut[17][5];
              muxOutConnector[49] = fifoOut[18][5];
              muxOutConnector[50] = fifoOut[19][5];
              muxOutConnector[51] = fifoOut[20][5];
       end
       7: begin
              muxOutConnector[0] = fifoOut[2][10];
              muxOutConnector[1] = fifoOut[3][10];
              muxOutConnector[2] = fifoOut[4][10];
              muxOutConnector[3] = fifoOut[5][10];
              muxOutConnector[4] = fifoOut[6][10];
              muxOutConnector[5] = fifoOut[7][10];
              muxOutConnector[6] = fifoOut[8][10];
              muxOutConnector[7] = fifoOut[9][10];
              muxOutConnector[8] = fifoOut[10][10];
              muxOutConnector[9] = fifoOut[11][10];
              muxOutConnector[10] = fifoOut[12][10];
              muxOutConnector[11] = fifoOut[13][10];
              muxOutConnector[12] = fifoOut[14][10];
              muxOutConnector[13] = fifoOut[15][10];
              muxOutConnector[14] = fifoOut[16][10];
              muxOutConnector[15] = fifoOut[17][10];
              muxOutConnector[16] = fifoOut[18][10];
              muxOutConnector[17] = fifoOut[19][10];
              muxOutConnector[18] = fifoOut[20][10];
              muxOutConnector[19] = fifoOut[21][10];
              muxOutConnector[20] = fifoOut[22][10];
              muxOutConnector[21] = fifoOut[23][10];
              muxOutConnector[22] = fifoOut[24][10];
              muxOutConnector[23] = fifoOut[25][10];
              muxOutConnector[24] = fifoOut[0][9];
              muxOutConnector[25] = fifoOut[1][9];
              muxOutConnector[26] = fifoOut[21][6];
              muxOutConnector[27] = fifoOut[22][6];
              muxOutConnector[28] = fifoOut[23][6];
              muxOutConnector[29] = fifoOut[24][6];
              muxOutConnector[30] = fifoOut[25][6];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = fifoOut[12][5];
              muxOutConnector[44] = fifoOut[13][5];
              muxOutConnector[45] = fifoOut[14][5];
              muxOutConnector[46] = fifoOut[15][5];
              muxOutConnector[47] = fifoOut[16][5];
              muxOutConnector[48] = fifoOut[17][5];
              muxOutConnector[49] = fifoOut[18][5];
              muxOutConnector[50] = fifoOut[19][5];
              muxOutConnector[51] = fifoOut[20][5];
       end
       8: begin
              muxOutConnector[0] = fifoOut[2][10];
              muxOutConnector[1] = fifoOut[3][10];
              muxOutConnector[2] = fifoOut[4][10];
              muxOutConnector[3] = fifoOut[5][10];
              muxOutConnector[4] = fifoOut[6][10];
              muxOutConnector[5] = fifoOut[7][10];
              muxOutConnector[6] = fifoOut[8][10];
              muxOutConnector[7] = fifoOut[9][10];
              muxOutConnector[8] = fifoOut[10][10];
              muxOutConnector[9] = fifoOut[11][10];
              muxOutConnector[10] = fifoOut[12][10];
              muxOutConnector[11] = fifoOut[13][10];
              muxOutConnector[12] = fifoOut[14][10];
              muxOutConnector[13] = fifoOut[15][10];
              muxOutConnector[14] = fifoOut[16][10];
              muxOutConnector[15] = fifoOut[17][10];
              muxOutConnector[16] = fifoOut[18][10];
              muxOutConnector[17] = fifoOut[19][10];
              muxOutConnector[18] = fifoOut[20][10];
              muxOutConnector[19] = fifoOut[21][10];
              muxOutConnector[20] = fifoOut[22][10];
              muxOutConnector[21] = fifoOut[23][10];
              muxOutConnector[22] = fifoOut[24][10];
              muxOutConnector[23] = fifoOut[25][10];
              muxOutConnector[24] = fifoOut[0][9];
              muxOutConnector[25] = fifoOut[1][9];
              muxOutConnector[26] = fifoOut[21][6];
              muxOutConnector[27] = fifoOut[22][6];
              muxOutConnector[28] = fifoOut[23][6];
              muxOutConnector[29] = fifoOut[24][6];
              muxOutConnector[30] = fifoOut[25][6];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = fifoOut[12][5];
              muxOutConnector[44] = fifoOut[13][5];
              muxOutConnector[45] = fifoOut[14][5];
              muxOutConnector[46] = fifoOut[15][5];
              muxOutConnector[47] = fifoOut[16][5];
              muxOutConnector[48] = fifoOut[17][5];
              muxOutConnector[49] = fifoOut[18][5];
              muxOutConnector[50] = fifoOut[19][5];
              muxOutConnector[51] = fifoOut[20][5];
       end
       9: begin
              muxOutConnector[0] = fifoOut[2][10];
              muxOutConnector[1] = fifoOut[3][10];
              muxOutConnector[2] = fifoOut[4][10];
              muxOutConnector[3] = fifoOut[5][10];
              muxOutConnector[4] = fifoOut[6][10];
              muxOutConnector[5] = fifoOut[7][10];
              muxOutConnector[6] = fifoOut[8][10];
              muxOutConnector[7] = fifoOut[9][10];
              muxOutConnector[8] = fifoOut[10][10];
              muxOutConnector[9] = fifoOut[11][10];
              muxOutConnector[10] = fifoOut[12][10];
              muxOutConnector[11] = fifoOut[13][10];
              muxOutConnector[12] = fifoOut[14][10];
              muxOutConnector[13] = fifoOut[15][10];
              muxOutConnector[14] = fifoOut[16][10];
              muxOutConnector[15] = fifoOut[17][10];
              muxOutConnector[16] = fifoOut[18][10];
              muxOutConnector[17] = fifoOut[19][10];
              muxOutConnector[18] = fifoOut[20][10];
              muxOutConnector[19] = fifoOut[21][10];
              muxOutConnector[20] = fifoOut[22][10];
              muxOutConnector[21] = fifoOut[23][10];
              muxOutConnector[22] = fifoOut[24][10];
              muxOutConnector[23] = fifoOut[25][10];
              muxOutConnector[24] = fifoOut[0][9];
              muxOutConnector[25] = fifoOut[1][9];
              muxOutConnector[26] = fifoOut[21][6];
              muxOutConnector[27] = fifoOut[22][6];
              muxOutConnector[28] = fifoOut[23][6];
              muxOutConnector[29] = fifoOut[24][6];
              muxOutConnector[30] = fifoOut[25][6];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = fifoOut[12][5];
              muxOutConnector[44] = fifoOut[13][5];
              muxOutConnector[45] = fifoOut[14][5];
              muxOutConnector[46] = fifoOut[15][5];
              muxOutConnector[47] = fifoOut[16][5];
              muxOutConnector[48] = fifoOut[17][5];
              muxOutConnector[49] = fifoOut[18][5];
              muxOutConnector[50] = fifoOut[19][5];
              muxOutConnector[51] = fifoOut[20][5];
       end
       10: begin
              muxOutConnector[0] = fifoOut[2][10];
              muxOutConnector[1] = fifoOut[3][10];
              muxOutConnector[2] = fifoOut[4][10];
              muxOutConnector[3] = fifoOut[5][10];
              muxOutConnector[4] = fifoOut[6][10];
              muxOutConnector[5] = fifoOut[7][10];
              muxOutConnector[6] = fifoOut[8][10];
              muxOutConnector[7] = fifoOut[9][10];
              muxOutConnector[8] = fifoOut[10][10];
              muxOutConnector[9] = fifoOut[11][10];
              muxOutConnector[10] = fifoOut[12][10];
              muxOutConnector[11] = fifoOut[13][10];
              muxOutConnector[12] = fifoOut[14][10];
              muxOutConnector[13] = fifoOut[15][10];
              muxOutConnector[14] = fifoOut[16][10];
              muxOutConnector[15] = fifoOut[26][9];
              muxOutConnector[16] = fifoOut[27][9];
              muxOutConnector[17] = fifoOut[28][9];
              muxOutConnector[18] = fifoOut[29][9];
              muxOutConnector[19] = fifoOut[30][9];
              muxOutConnector[20] = fifoOut[31][9];
              muxOutConnector[21] = fifoOut[32][9];
              muxOutConnector[22] = fifoOut[33][9];
              muxOutConnector[23] = fifoOut[34][9];
              muxOutConnector[24] = fifoOut[35][9];
              muxOutConnector[25] = fifoOut[36][9];
              muxOutConnector[26] = fifoOut[21][6];
              muxOutConnector[27] = fifoOut[22][6];
              muxOutConnector[28] = fifoOut[23][6];
              muxOutConnector[29] = fifoOut[24][6];
              muxOutConnector[30] = fifoOut[25][6];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = fifoOut[12][5];
              muxOutConnector[44] = fifoOut[13][5];
              muxOutConnector[45] = fifoOut[14][5];
              muxOutConnector[46] = fifoOut[15][5];
              muxOutConnector[47] = fifoOut[16][5];
              muxOutConnector[48] = fifoOut[17][5];
              muxOutConnector[49] = fifoOut[18][5];
              muxOutConnector[50] = fifoOut[19][5];
              muxOutConnector[51] = fifoOut[20][5];
       end
       11: begin
              muxOutConnector[0] = fifoOut[37][10];
              muxOutConnector[1] = fifoOut[38][10];
              muxOutConnector[2] = fifoOut[39][10];
              muxOutConnector[3] = fifoOut[40][10];
              muxOutConnector[4] = fifoOut[41][10];
              muxOutConnector[5] = fifoOut[42][10];
              muxOutConnector[6] = fifoOut[43][10];
              muxOutConnector[7] = fifoOut[44][10];
              muxOutConnector[8] = fifoOut[45][10];
              muxOutConnector[9] = fifoOut[46][10];
              muxOutConnector[10] = fifoOut[47][10];
              muxOutConnector[11] = fifoOut[48][10];
              muxOutConnector[12] = fifoOut[49][10];
              muxOutConnector[13] = fifoOut[50][10];
              muxOutConnector[14] = fifoOut[51][10];
              muxOutConnector[15] = fifoOut[26][9];
              muxOutConnector[16] = fifoOut[27][9];
              muxOutConnector[17] = fifoOut[28][9];
              muxOutConnector[18] = fifoOut[29][9];
              muxOutConnector[19] = fifoOut[30][9];
              muxOutConnector[20] = fifoOut[31][9];
              muxOutConnector[21] = fifoOut[32][9];
              muxOutConnector[22] = fifoOut[33][9];
              muxOutConnector[23] = fifoOut[34][9];
              muxOutConnector[24] = fifoOut[35][9];
              muxOutConnector[25] = fifoOut[36][9];
              muxOutConnector[26] = fifoOut[21][6];
              muxOutConnector[27] = fifoOut[22][6];
              muxOutConnector[28] = fifoOut[23][6];
              muxOutConnector[29] = fifoOut[24][6];
              muxOutConnector[30] = fifoOut[25][6];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = fifoOut[12][5];
              muxOutConnector[44] = fifoOut[13][5];
              muxOutConnector[45] = fifoOut[14][5];
              muxOutConnector[46] = fifoOut[15][5];
              muxOutConnector[47] = fifoOut[16][5];
              muxOutConnector[48] = fifoOut[17][5];
              muxOutConnector[49] = fifoOut[18][5];
              muxOutConnector[50] = fifoOut[19][5];
              muxOutConnector[51] = fifoOut[20][5];
       end
       12: begin
              muxOutConnector[0] = fifoOut[37][10];
              muxOutConnector[1] = fifoOut[38][10];
              muxOutConnector[2] = fifoOut[39][10];
              muxOutConnector[3] = fifoOut[40][10];
              muxOutConnector[4] = fifoOut[41][10];
              muxOutConnector[5] = fifoOut[42][10];
              muxOutConnector[6] = fifoOut[43][10];
              muxOutConnector[7] = fifoOut[44][10];
              muxOutConnector[8] = fifoOut[45][10];
              muxOutConnector[9] = fifoOut[46][10];
              muxOutConnector[10] = fifoOut[47][10];
              muxOutConnector[11] = fifoOut[48][10];
              muxOutConnector[12] = fifoOut[49][10];
              muxOutConnector[13] = fifoOut[50][10];
              muxOutConnector[14] = fifoOut[51][10];
              muxOutConnector[15] = fifoOut[26][9];
              muxOutConnector[16] = fifoOut[27][9];
              muxOutConnector[17] = fifoOut[28][9];
              muxOutConnector[18] = fifoOut[29][9];
              muxOutConnector[19] = fifoOut[30][9];
              muxOutConnector[20] = fifoOut[31][9];
              muxOutConnector[21] = fifoOut[32][9];
              muxOutConnector[22] = fifoOut[33][9];
              muxOutConnector[23] = fifoOut[34][9];
              muxOutConnector[24] = fifoOut[35][9];
              muxOutConnector[25] = fifoOut[36][9];
              muxOutConnector[26] = fifoOut[21][6];
              muxOutConnector[27] = fifoOut[22][6];
              muxOutConnector[28] = fifoOut[23][6];
              muxOutConnector[29] = fifoOut[24][6];
              muxOutConnector[30] = fifoOut[25][6];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = fifoOut[12][5];
              muxOutConnector[44] = fifoOut[13][5];
              muxOutConnector[45] = fifoOut[14][5];
              muxOutConnector[46] = fifoOut[15][5];
              muxOutConnector[47] = fifoOut[16][5];
              muxOutConnector[48] = fifoOut[17][5];
              muxOutConnector[49] = fifoOut[18][5];
              muxOutConnector[50] = fifoOut[19][5];
              muxOutConnector[51] = fifoOut[20][5];
       end
       13: begin
              muxOutConnector[0] = fifoOut[37][10];
              muxOutConnector[1] = fifoOut[38][10];
              muxOutConnector[2] = fifoOut[39][10];
              muxOutConnector[3] = fifoOut[40][10];
              muxOutConnector[4] = fifoOut[41][10];
              muxOutConnector[5] = fifoOut[42][10];
              muxOutConnector[6] = fifoOut[43][10];
              muxOutConnector[7] = fifoOut[44][10];
              muxOutConnector[8] = fifoOut[45][10];
              muxOutConnector[9] = fifoOut[46][10];
              muxOutConnector[10] = fifoOut[47][10];
              muxOutConnector[11] = fifoOut[48][10];
              muxOutConnector[12] = fifoOut[49][10];
              muxOutConnector[13] = fifoOut[50][10];
              muxOutConnector[14] = fifoOut[51][10];
              muxOutConnector[15] = fifoOut[26][9];
              muxOutConnector[16] = fifoOut[27][9];
              muxOutConnector[17] = fifoOut[28][9];
              muxOutConnector[18] = fifoOut[29][9];
              muxOutConnector[19] = fifoOut[30][9];
              muxOutConnector[20] = fifoOut[31][9];
              muxOutConnector[21] = fifoOut[32][9];
              muxOutConnector[22] = fifoOut[33][9];
              muxOutConnector[23] = fifoOut[34][9];
              muxOutConnector[24] = fifoOut[35][9];
              muxOutConnector[25] = fifoOut[36][9];
              muxOutConnector[26] = fifoOut[21][6];
              muxOutConnector[27] = fifoOut[22][6];
              muxOutConnector[28] = fifoOut[23][6];
              muxOutConnector[29] = fifoOut[24][6];
              muxOutConnector[30] = fifoOut[25][6];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = fifoOut[12][5];
              muxOutConnector[44] = fifoOut[13][5];
              muxOutConnector[45] = fifoOut[14][5];
              muxOutConnector[46] = fifoOut[15][5];
              muxOutConnector[47] = fifoOut[16][5];
              muxOutConnector[48] = fifoOut[17][5];
              muxOutConnector[49] = fifoOut[18][5];
              muxOutConnector[50] = fifoOut[19][5];
              muxOutConnector[51] = fifoOut[20][5];
       end
       14: begin
              muxOutConnector[0] = fifoOut[37][10];
              muxOutConnector[1] = fifoOut[38][10];
              muxOutConnector[2] = fifoOut[39][10];
              muxOutConnector[3] = fifoOut[40][10];
              muxOutConnector[4] = fifoOut[41][10];
              muxOutConnector[5] = fifoOut[42][10];
              muxOutConnector[6] = fifoOut[43][10];
              muxOutConnector[7] = fifoOut[44][10];
              muxOutConnector[8] = fifoOut[45][10];
              muxOutConnector[9] = fifoOut[46][10];
              muxOutConnector[10] = fifoOut[47][10];
              muxOutConnector[11] = fifoOut[48][10];
              muxOutConnector[12] = fifoOut[49][10];
              muxOutConnector[13] = fifoOut[50][10];
              muxOutConnector[14] = fifoOut[51][10];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[2][13];
              muxOutConnector[18] = fifoOut[3][13];
              muxOutConnector[19] = fifoOut[4][13];
              muxOutConnector[20] = fifoOut[5][13];
              muxOutConnector[21] = fifoOut[6][13];
              muxOutConnector[22] = fifoOut[7][13];
              muxOutConnector[23] = fifoOut[8][13];
              muxOutConnector[24] = fifoOut[9][13];
              muxOutConnector[25] = fifoOut[10][13];
              muxOutConnector[26] = fifoOut[21][6];
              muxOutConnector[27] = fifoOut[22][6];
              muxOutConnector[28] = fifoOut[23][6];
              muxOutConnector[29] = fifoOut[24][6];
              muxOutConnector[30] = fifoOut[25][6];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = fifoOut[12][5];
              muxOutConnector[44] = fifoOut[13][5];
              muxOutConnector[45] = fifoOut[14][5];
              muxOutConnector[46] = fifoOut[15][5];
              muxOutConnector[47] = fifoOut[16][5];
              muxOutConnector[48] = fifoOut[17][5];
              muxOutConnector[49] = fifoOut[18][5];
              muxOutConnector[50] = fifoOut[19][5];
              muxOutConnector[51] = fifoOut[20][5];
       end
       15: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[2][13];
              muxOutConnector[18] = fifoOut[3][13];
              muxOutConnector[19] = fifoOut[4][13];
              muxOutConnector[20] = fifoOut[5][13];
              muxOutConnector[21] = fifoOut[6][13];
              muxOutConnector[22] = fifoOut[7][13];
              muxOutConnector[23] = fifoOut[8][13];
              muxOutConnector[24] = fifoOut[9][13];
              muxOutConnector[25] = fifoOut[10][13];
              muxOutConnector[26] = fifoOut[21][6];
              muxOutConnector[27] = fifoOut[22][6];
              muxOutConnector[28] = fifoOut[23][6];
              muxOutConnector[29] = fifoOut[24][6];
              muxOutConnector[30] = fifoOut[25][6];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = fifoOut[12][5];
              muxOutConnector[44] = fifoOut[13][5];
              muxOutConnector[45] = fifoOut[14][5];
              muxOutConnector[46] = fifoOut[15][5];
              muxOutConnector[47] = fifoOut[16][5];
              muxOutConnector[48] = fifoOut[17][5];
              muxOutConnector[49] = fifoOut[18][5];
              muxOutConnector[50] = fifoOut[19][5];
              muxOutConnector[51] = fifoOut[20][5];
       end
       16: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[2][13];
              muxOutConnector[18] = fifoOut[3][13];
              muxOutConnector[19] = fifoOut[4][13];
              muxOutConnector[20] = fifoOut[5][13];
              muxOutConnector[21] = fifoOut[6][13];
              muxOutConnector[22] = fifoOut[7][13];
              muxOutConnector[23] = fifoOut[8][13];
              muxOutConnector[24] = fifoOut[9][13];
              muxOutConnector[25] = fifoOut[10][13];
              muxOutConnector[26] = fifoOut[21][6];
              muxOutConnector[27] = fifoOut[22][6];
              muxOutConnector[28] = fifoOut[23][6];
              muxOutConnector[29] = fifoOut[24][6];
              muxOutConnector[30] = fifoOut[25][6];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = fifoOut[12][5];
              muxOutConnector[44] = fifoOut[13][5];
              muxOutConnector[45] = fifoOut[14][5];
              muxOutConnector[46] = fifoOut[15][5];
              muxOutConnector[47] = fifoOut[16][5];
              muxOutConnector[48] = fifoOut[17][5];
              muxOutConnector[49] = fifoOut[18][5];
              muxOutConnector[50] = fifoOut[19][5];
              muxOutConnector[51] = fifoOut[20][5];
       end
       17: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[2][13];
              muxOutConnector[18] = fifoOut[3][13];
              muxOutConnector[19] = fifoOut[4][13];
              muxOutConnector[20] = fifoOut[5][13];
              muxOutConnector[21] = fifoOut[6][13];
              muxOutConnector[22] = fifoOut[7][13];
              muxOutConnector[23] = fifoOut[8][13];
              muxOutConnector[24] = fifoOut[9][13];
              muxOutConnector[25] = fifoOut[10][13];
              muxOutConnector[26] = fifoOut[21][6];
              muxOutConnector[27] = fifoOut[22][6];
              muxOutConnector[28] = fifoOut[23][6];
              muxOutConnector[29] = fifoOut[24][6];
              muxOutConnector[30] = fifoOut[25][6];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = fifoOut[12][5];
              muxOutConnector[44] = fifoOut[13][5];
              muxOutConnector[45] = fifoOut[14][5];
              muxOutConnector[46] = fifoOut[15][5];
              muxOutConnector[47] = fifoOut[16][5];
              muxOutConnector[48] = fifoOut[17][5];
              muxOutConnector[49] = fifoOut[18][5];
              muxOutConnector[50] = fifoOut[19][5];
              muxOutConnector[51] = fifoOut[20][5];
       end
       18: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[2][13];
              muxOutConnector[18] = fifoOut[3][13];
              muxOutConnector[19] = fifoOut[4][13];
              muxOutConnector[20] = fifoOut[5][13];
              muxOutConnector[21] = fifoOut[6][13];
              muxOutConnector[22] = fifoOut[7][13];
              muxOutConnector[23] = fifoOut[8][13];
              muxOutConnector[24] = fifoOut[9][13];
              muxOutConnector[25] = fifoOut[10][13];
              muxOutConnector[26] = fifoOut[21][6];
              muxOutConnector[27] = fifoOut[22][6];
              muxOutConnector[28] = fifoOut[23][6];
              muxOutConnector[29] = fifoOut[24][6];
              muxOutConnector[30] = fifoOut[25][6];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = fifoOut[12][5];
              muxOutConnector[44] = fifoOut[13][5];
              muxOutConnector[45] = fifoOut[14][5];
              muxOutConnector[46] = fifoOut[15][5];
              muxOutConnector[47] = fifoOut[16][5];
              muxOutConnector[48] = fifoOut[17][5];
              muxOutConnector[49] = fifoOut[18][5];
              muxOutConnector[50] = fifoOut[19][5];
              muxOutConnector[51] = fifoOut[20][5];
       end
       19: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[21][6];
              muxOutConnector[27] = fifoOut[22][6];
              muxOutConnector[28] = fifoOut[23][6];
              muxOutConnector[29] = fifoOut[24][6];
              muxOutConnector[30] = fifoOut[25][6];
              muxOutConnector[31] = fifoOut[0][5];
              muxOutConnector[32] = fifoOut[1][5];
              muxOutConnector[33] = fifoOut[2][5];
              muxOutConnector[34] = fifoOut[3][5];
              muxOutConnector[35] = fifoOut[4][5];
              muxOutConnector[36] = fifoOut[5][5];
              muxOutConnector[37] = fifoOut[6][5];
              muxOutConnector[38] = fifoOut[7][5];
              muxOutConnector[39] = fifoOut[8][5];
              muxOutConnector[40] = fifoOut[9][5];
              muxOutConnector[41] = fifoOut[10][5];
              muxOutConnector[42] = fifoOut[11][5];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
