`timescale 1ns / 1ps
module LMem1To0_511_circ4_combined_ys_yu_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        rxIn,
        load_input_en,
        iteration_0_indicator,
        feedback_en,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter r_lower = 32;
parameter c = 17;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input load_input_en;
input iteration_0_indicator;
input [ADDRESSWIDTH-1:0]unloadAddress;
input feedback_en;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input [ r_lower * w - 1 : 0 ] rxIn; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
wire [w-1:0]rxInConnector[r_lower-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

generate
    for (k=0;k<r_lower;k=k+1)begin:assign_rx
        assign rxInConnector[k] = rxIn[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            if(feedback_en)begin
                 fifoOut[i][0] <= fifoOut[i][c-1];
            end
            else if(load_input_en)begin
                 if(i < r_lower)begin
                   fifoOut[i][0] = rxInConnector[i];
                 end
                 else begin
                   fifoOut[i][0] = maxVal;
                 end
            end
            else begin
                 fifoOut[i][0] <= ly0InConnector[i];
            end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
       0: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = fifoOut[10][8][w-1];
              unloadMuxOut[29] = fifoOut[11][8][w-1];
              unloadMuxOut[30] = fifoOut[12][8][w-1];
              unloadMuxOut[31] = fifoOut[13][8][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[14][9][w-1];
              unloadMuxOut[1] = fifoOut[15][9][w-1];
              unloadMuxOut[2] = fifoOut[16][9][w-1];
              unloadMuxOut[3] = fifoOut[17][9][w-1];
              unloadMuxOut[4] = fifoOut[18][9][w-1];
              unloadMuxOut[5] = fifoOut[19][9][w-1];
              unloadMuxOut[6] = fifoOut[20][9][w-1];
              unloadMuxOut[7] = fifoOut[21][9][w-1];
              unloadMuxOut[8] = fifoOut[22][9][w-1];
              unloadMuxOut[9] = fifoOut[23][9][w-1];
              unloadMuxOut[10] = fifoOut[24][9][w-1];
              unloadMuxOut[11] = fifoOut[25][9][w-1];
              unloadMuxOut[12] = fifoOut[0][8][w-1];
              unloadMuxOut[13] = fifoOut[1][8][w-1];
              unloadMuxOut[14] = fifoOut[2][8][w-1];
              unloadMuxOut[15] = fifoOut[3][8][w-1];
              unloadMuxOut[16] = fifoOut[4][8][w-1];
              unloadMuxOut[17] = fifoOut[5][8][w-1];
              unloadMuxOut[18] = fifoOut[6][8][w-1];
              unloadMuxOut[19] = fifoOut[7][8][w-1];
              unloadMuxOut[20] = fifoOut[8][8][w-1];
              unloadMuxOut[21] = fifoOut[9][8][w-1];
              unloadMuxOut[22] = fifoOut[10][8][w-1];
              unloadMuxOut[23] = fifoOut[11][8][w-1];
              unloadMuxOut[24] = fifoOut[12][8][w-1];
              unloadMuxOut[25] = fifoOut[13][8][w-1];
              unloadMuxOut[26] = fifoOut[14][8][w-1];
              unloadMuxOut[27] = fifoOut[15][8][w-1];
              unloadMuxOut[28] = fifoOut[16][8][w-1];
              unloadMuxOut[29] = fifoOut[17][8][w-1];
              unloadMuxOut[30] = fifoOut[18][8][w-1];
              unloadMuxOut[31] = fifoOut[19][8][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[20][9][w-1];
              unloadMuxOut[1] = fifoOut[21][9][w-1];
              unloadMuxOut[2] = fifoOut[22][9][w-1];
              unloadMuxOut[3] = fifoOut[23][9][w-1];
              unloadMuxOut[4] = fifoOut[24][9][w-1];
              unloadMuxOut[5] = fifoOut[25][9][w-1];
              unloadMuxOut[6] = fifoOut[0][8][w-1];
              unloadMuxOut[7] = fifoOut[1][8][w-1];
              unloadMuxOut[8] = fifoOut[2][8][w-1];
              unloadMuxOut[9] = fifoOut[3][8][w-1];
              unloadMuxOut[10] = fifoOut[4][8][w-1];
              unloadMuxOut[11] = fifoOut[5][8][w-1];
              unloadMuxOut[12] = fifoOut[6][8][w-1];
              unloadMuxOut[13] = fifoOut[7][8][w-1];
              unloadMuxOut[14] = fifoOut[8][8][w-1];
              unloadMuxOut[15] = fifoOut[9][8][w-1];
              unloadMuxOut[16] = fifoOut[10][8][w-1];
              unloadMuxOut[17] = fifoOut[11][8][w-1];
              unloadMuxOut[18] = fifoOut[12][8][w-1];
              unloadMuxOut[19] = fifoOut[13][8][w-1];
              unloadMuxOut[20] = fifoOut[14][8][w-1];
              unloadMuxOut[21] = fifoOut[15][8][w-1];
              unloadMuxOut[22] = fifoOut[16][8][w-1];
              unloadMuxOut[23] = fifoOut[17][8][w-1];
              unloadMuxOut[24] = fifoOut[18][8][w-1];
              unloadMuxOut[25] = fifoOut[19][8][w-1];
              unloadMuxOut[26] = fifoOut[20][8][w-1];
              unloadMuxOut[27] = fifoOut[21][8][w-1];
              unloadMuxOut[28] = fifoOut[22][8][w-1];
              unloadMuxOut[29] = fifoOut[23][8][w-1];
              unloadMuxOut[30] = fifoOut[24][8][w-1];
              unloadMuxOut[31] = fifoOut[25][8][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[0][8][w-1];
              unloadMuxOut[1] = fifoOut[1][8][w-1];
              unloadMuxOut[2] = fifoOut[2][8][w-1];
              unloadMuxOut[3] = fifoOut[3][8][w-1];
              unloadMuxOut[4] = fifoOut[4][8][w-1];
              unloadMuxOut[5] = fifoOut[5][8][w-1];
              unloadMuxOut[6] = fifoOut[6][8][w-1];
              unloadMuxOut[7] = fifoOut[7][8][w-1];
              unloadMuxOut[8] = fifoOut[8][8][w-1];
              unloadMuxOut[9] = fifoOut[9][8][w-1];
              unloadMuxOut[10] = fifoOut[10][8][w-1];
              unloadMuxOut[11] = fifoOut[11][8][w-1];
              unloadMuxOut[12] = fifoOut[12][8][w-1];
              unloadMuxOut[13] = fifoOut[13][8][w-1];
              unloadMuxOut[14] = fifoOut[14][8][w-1];
              unloadMuxOut[15] = fifoOut[15][8][w-1];
              unloadMuxOut[16] = fifoOut[16][8][w-1];
              unloadMuxOut[17] = fifoOut[17][8][w-1];
              unloadMuxOut[18] = fifoOut[18][8][w-1];
              unloadMuxOut[19] = fifoOut[19][8][w-1];
              unloadMuxOut[20] = fifoOut[20][8][w-1];
              unloadMuxOut[21] = fifoOut[21][8][w-1];
              unloadMuxOut[22] = fifoOut[22][8][w-1];
              unloadMuxOut[23] = fifoOut[26][15][w-1];
              unloadMuxOut[24] = fifoOut[27][15][w-1];
              unloadMuxOut[25] = fifoOut[28][15][w-1];
              unloadMuxOut[26] = fifoOut[29][15][w-1];
              unloadMuxOut[27] = fifoOut[30][15][w-1];
              unloadMuxOut[28] = fifoOut[31][15][w-1];
              unloadMuxOut[29] = fifoOut[32][15][w-1];
              unloadMuxOut[30] = fifoOut[33][15][w-1];
              unloadMuxOut[31] = fifoOut[34][15][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[35][16][w-1];
              unloadMuxOut[1] = fifoOut[36][16][w-1];
              unloadMuxOut[2] = fifoOut[37][16][w-1];
              unloadMuxOut[3] = fifoOut[38][16][w-1];
              unloadMuxOut[4] = fifoOut[39][16][w-1];
              unloadMuxOut[5] = fifoOut[40][16][w-1];
              unloadMuxOut[6] = fifoOut[41][16][w-1];
              unloadMuxOut[7] = fifoOut[42][16][w-1];
              unloadMuxOut[8] = fifoOut[43][16][w-1];
              unloadMuxOut[9] = fifoOut[44][16][w-1];
              unloadMuxOut[10] = fifoOut[45][16][w-1];
              unloadMuxOut[11] = fifoOut[46][16][w-1];
              unloadMuxOut[12] = fifoOut[47][16][w-1];
              unloadMuxOut[13] = fifoOut[48][16][w-1];
              unloadMuxOut[14] = fifoOut[49][16][w-1];
              unloadMuxOut[15] = fifoOut[50][16][w-1];
              unloadMuxOut[16] = fifoOut[51][16][w-1];
              unloadMuxOut[17] = fifoOut[26][15][w-1];
              unloadMuxOut[18] = fifoOut[27][15][w-1];
              unloadMuxOut[19] = fifoOut[28][15][w-1];
              unloadMuxOut[20] = fifoOut[29][15][w-1];
              unloadMuxOut[21] = fifoOut[30][15][w-1];
              unloadMuxOut[22] = fifoOut[31][15][w-1];
              unloadMuxOut[23] = fifoOut[32][15][w-1];
              unloadMuxOut[24] = fifoOut[33][15][w-1];
              unloadMuxOut[25] = fifoOut[34][15][w-1];
              unloadMuxOut[26] = fifoOut[35][15][w-1];
              unloadMuxOut[27] = fifoOut[36][15][w-1];
              unloadMuxOut[28] = fifoOut[37][15][w-1];
              unloadMuxOut[29] = fifoOut[38][15][w-1];
              unloadMuxOut[30] = fifoOut[39][15][w-1];
              unloadMuxOut[31] = fifoOut[40][15][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[41][16][w-1];
              unloadMuxOut[1] = fifoOut[42][16][w-1];
              unloadMuxOut[2] = fifoOut[43][16][w-1];
              unloadMuxOut[3] = fifoOut[44][16][w-1];
              unloadMuxOut[4] = fifoOut[45][16][w-1];
              unloadMuxOut[5] = fifoOut[46][16][w-1];
              unloadMuxOut[6] = fifoOut[47][16][w-1];
              unloadMuxOut[7] = fifoOut[48][16][w-1];
              unloadMuxOut[8] = fifoOut[49][16][w-1];
              unloadMuxOut[9] = fifoOut[50][16][w-1];
              unloadMuxOut[10] = fifoOut[51][16][w-1];
              unloadMuxOut[11] = fifoOut[26][15][w-1];
              unloadMuxOut[12] = fifoOut[27][15][w-1];
              unloadMuxOut[13] = fifoOut[28][15][w-1];
              unloadMuxOut[14] = fifoOut[29][15][w-1];
              unloadMuxOut[15] = fifoOut[30][15][w-1];
              unloadMuxOut[16] = fifoOut[31][15][w-1];
              unloadMuxOut[17] = fifoOut[32][15][w-1];
              unloadMuxOut[18] = fifoOut[33][15][w-1];
              unloadMuxOut[19] = fifoOut[34][15][w-1];
              unloadMuxOut[20] = fifoOut[35][15][w-1];
              unloadMuxOut[21] = fifoOut[36][15][w-1];
              unloadMuxOut[22] = fifoOut[37][15][w-1];
              unloadMuxOut[23] = fifoOut[38][15][w-1];
              unloadMuxOut[24] = fifoOut[39][15][w-1];
              unloadMuxOut[25] = fifoOut[40][15][w-1];
              unloadMuxOut[26] = fifoOut[41][15][w-1];
              unloadMuxOut[27] = fifoOut[42][15][w-1];
              unloadMuxOut[28] = fifoOut[43][15][w-1];
              unloadMuxOut[29] = fifoOut[44][15][w-1];
              unloadMuxOut[30] = fifoOut[45][15][w-1];
              unloadMuxOut[31] = fifoOut[46][15][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[47][16][w-1];
              unloadMuxOut[1] = fifoOut[48][16][w-1];
              unloadMuxOut[2] = fifoOut[49][16][w-1];
              unloadMuxOut[3] = fifoOut[50][16][w-1];
              unloadMuxOut[4] = fifoOut[51][16][w-1];
              unloadMuxOut[5] = fifoOut[26][15][w-1];
              unloadMuxOut[6] = fifoOut[27][15][w-1];
              unloadMuxOut[7] = fifoOut[28][15][w-1];
              unloadMuxOut[8] = fifoOut[29][15][w-1];
              unloadMuxOut[9] = fifoOut[30][15][w-1];
              unloadMuxOut[10] = fifoOut[31][15][w-1];
              unloadMuxOut[11] = fifoOut[32][15][w-1];
              unloadMuxOut[12] = fifoOut[33][15][w-1];
              unloadMuxOut[13] = fifoOut[34][15][w-1];
              unloadMuxOut[14] = fifoOut[35][15][w-1];
              unloadMuxOut[15] = fifoOut[36][15][w-1];
              unloadMuxOut[16] = fifoOut[37][15][w-1];
              unloadMuxOut[17] = fifoOut[38][15][w-1];
              unloadMuxOut[18] = fifoOut[39][15][w-1];
              unloadMuxOut[19] = fifoOut[40][15][w-1];
              unloadMuxOut[20] = fifoOut[41][15][w-1];
              unloadMuxOut[21] = fifoOut[42][15][w-1];
              unloadMuxOut[22] = fifoOut[43][15][w-1];
              unloadMuxOut[23] = fifoOut[44][15][w-1];
              unloadMuxOut[24] = fifoOut[45][15][w-1];
              unloadMuxOut[25] = fifoOut[46][15][w-1];
              unloadMuxOut[26] = fifoOut[47][15][w-1];
              unloadMuxOut[27] = fifoOut[48][15][w-1];
              unloadMuxOut[28] = fifoOut[49][15][w-1];
              unloadMuxOut[29] = fifoOut[50][15][w-1];
              unloadMuxOut[30] = fifoOut[51][15][w-1];
              unloadMuxOut[31] = fifoOut[26][14][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[27][15][w-1];
              unloadMuxOut[1] = fifoOut[28][15][w-1];
              unloadMuxOut[2] = fifoOut[29][15][w-1];
              unloadMuxOut[3] = fifoOut[30][15][w-1];
              unloadMuxOut[4] = fifoOut[31][15][w-1];
              unloadMuxOut[5] = fifoOut[32][15][w-1];
              unloadMuxOut[6] = fifoOut[33][15][w-1];
              unloadMuxOut[7] = fifoOut[34][15][w-1];
              unloadMuxOut[8] = fifoOut[35][15][w-1];
              unloadMuxOut[9] = fifoOut[36][15][w-1];
              unloadMuxOut[10] = fifoOut[37][15][w-1];
              unloadMuxOut[11] = fifoOut[38][15][w-1];
              unloadMuxOut[12] = fifoOut[39][15][w-1];
              unloadMuxOut[13] = fifoOut[40][15][w-1];
              unloadMuxOut[14] = fifoOut[41][15][w-1];
              unloadMuxOut[15] = fifoOut[42][15][w-1];
              unloadMuxOut[16] = fifoOut[43][15][w-1];
              unloadMuxOut[17] = fifoOut[44][15][w-1];
              unloadMuxOut[18] = fifoOut[45][15][w-1];
              unloadMuxOut[19] = fifoOut[46][15][w-1];
              unloadMuxOut[20] = fifoOut[47][15][w-1];
              unloadMuxOut[21] = fifoOut[48][15][w-1];
              unloadMuxOut[22] = fifoOut[49][15][w-1];
              unloadMuxOut[23] = fifoOut[50][15][w-1];
              unloadMuxOut[24] = fifoOut[51][15][w-1];
              unloadMuxOut[25] = fifoOut[26][14][w-1];
              unloadMuxOut[26] = fifoOut[27][14][w-1];
              unloadMuxOut[27] = fifoOut[28][14][w-1];
              unloadMuxOut[28] = fifoOut[29][14][w-1];
              unloadMuxOut[29] = fifoOut[30][14][w-1];
              unloadMuxOut[30] = fifoOut[31][14][w-1];
              unloadMuxOut[31] = fifoOut[32][14][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[33][15][w-1];
              unloadMuxOut[1] = fifoOut[34][15][w-1];
              unloadMuxOut[2] = fifoOut[35][15][w-1];
              unloadMuxOut[3] = fifoOut[36][15][w-1];
              unloadMuxOut[4] = fifoOut[37][15][w-1];
              unloadMuxOut[5] = fifoOut[38][15][w-1];
              unloadMuxOut[6] = fifoOut[39][15][w-1];
              unloadMuxOut[7] = fifoOut[40][15][w-1];
              unloadMuxOut[8] = fifoOut[41][15][w-1];
              unloadMuxOut[9] = fifoOut[42][15][w-1];
              unloadMuxOut[10] = fifoOut[43][15][w-1];
              unloadMuxOut[11] = fifoOut[44][15][w-1];
              unloadMuxOut[12] = fifoOut[45][15][w-1];
              unloadMuxOut[13] = fifoOut[46][15][w-1];
              unloadMuxOut[14] = fifoOut[47][15][w-1];
              unloadMuxOut[15] = fifoOut[48][15][w-1];
              unloadMuxOut[16] = fifoOut[49][15][w-1];
              unloadMuxOut[17] = fifoOut[50][15][w-1];
              unloadMuxOut[18] = fifoOut[51][15][w-1];
              unloadMuxOut[19] = fifoOut[26][14][w-1];
              unloadMuxOut[20] = fifoOut[27][14][w-1];
              unloadMuxOut[21] = fifoOut[28][14][w-1];
              unloadMuxOut[22] = fifoOut[29][14][w-1];
              unloadMuxOut[23] = fifoOut[30][14][w-1];
              unloadMuxOut[24] = fifoOut[31][14][w-1];
              unloadMuxOut[25] = fifoOut[32][14][w-1];
              unloadMuxOut[26] = fifoOut[33][14][w-1];
              unloadMuxOut[27] = fifoOut[34][14][w-1];
              unloadMuxOut[28] = fifoOut[35][14][w-1];
              unloadMuxOut[29] = fifoOut[36][14][w-1];
              unloadMuxOut[30] = fifoOut[37][14][w-1];
              unloadMuxOut[31] = fifoOut[38][14][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[39][15][w-1];
              unloadMuxOut[1] = fifoOut[40][15][w-1];
              unloadMuxOut[2] = fifoOut[41][15][w-1];
              unloadMuxOut[3] = fifoOut[42][15][w-1];
              unloadMuxOut[4] = fifoOut[43][15][w-1];
              unloadMuxOut[5] = fifoOut[44][15][w-1];
              unloadMuxOut[6] = fifoOut[45][15][w-1];
              unloadMuxOut[7] = fifoOut[46][15][w-1];
              unloadMuxOut[8] = fifoOut[47][15][w-1];
              unloadMuxOut[9] = fifoOut[48][15][w-1];
              unloadMuxOut[10] = fifoOut[49][15][w-1];
              unloadMuxOut[11] = fifoOut[50][15][w-1];
              unloadMuxOut[12] = fifoOut[51][15][w-1];
              unloadMuxOut[13] = fifoOut[26][14][w-1];
              unloadMuxOut[14] = fifoOut[27][14][w-1];
              unloadMuxOut[15] = fifoOut[28][14][w-1];
              unloadMuxOut[16] = fifoOut[29][14][w-1];
              unloadMuxOut[17] = fifoOut[30][14][w-1];
              unloadMuxOut[18] = fifoOut[31][14][w-1];
              unloadMuxOut[19] = fifoOut[32][14][w-1];
              unloadMuxOut[20] = fifoOut[33][14][w-1];
              unloadMuxOut[21] = fifoOut[34][14][w-1];
              unloadMuxOut[22] = fifoOut[35][14][w-1];
              unloadMuxOut[23] = fifoOut[36][14][w-1];
              unloadMuxOut[24] = fifoOut[37][14][w-1];
              unloadMuxOut[25] = fifoOut[38][14][w-1];
              unloadMuxOut[26] = fifoOut[39][14][w-1];
              unloadMuxOut[27] = fifoOut[40][14][w-1];
              unloadMuxOut[28] = fifoOut[41][14][w-1];
              unloadMuxOut[29] = fifoOut[42][14][w-1];
              unloadMuxOut[30] = fifoOut[43][14][w-1];
              unloadMuxOut[31] = fifoOut[44][14][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[45][15][w-1];
              unloadMuxOut[1] = fifoOut[46][15][w-1];
              unloadMuxOut[2] = fifoOut[47][15][w-1];
              unloadMuxOut[3] = fifoOut[48][15][w-1];
              unloadMuxOut[4] = fifoOut[49][15][w-1];
              unloadMuxOut[5] = fifoOut[50][15][w-1];
              unloadMuxOut[6] = fifoOut[51][15][w-1];
              unloadMuxOut[7] = fifoOut[26][14][w-1];
              unloadMuxOut[8] = fifoOut[27][14][w-1];
              unloadMuxOut[9] = fifoOut[28][14][w-1];
              unloadMuxOut[10] = fifoOut[29][14][w-1];
              unloadMuxOut[11] = fifoOut[30][14][w-1];
              unloadMuxOut[12] = fifoOut[31][14][w-1];
              unloadMuxOut[13] = fifoOut[32][14][w-1];
              unloadMuxOut[14] = fifoOut[33][14][w-1];
              unloadMuxOut[15] = fifoOut[34][14][w-1];
              unloadMuxOut[16] = fifoOut[35][14][w-1];
              unloadMuxOut[17] = fifoOut[36][14][w-1];
              unloadMuxOut[18] = fifoOut[37][14][w-1];
              unloadMuxOut[19] = fifoOut[38][14][w-1];
              unloadMuxOut[20] = fifoOut[39][14][w-1];
              unloadMuxOut[21] = fifoOut[40][14][w-1];
              unloadMuxOut[22] = fifoOut[41][14][w-1];
              unloadMuxOut[23] = fifoOut[42][14][w-1];
              unloadMuxOut[24] = fifoOut[43][14][w-1];
              unloadMuxOut[25] = fifoOut[44][14][w-1];
              unloadMuxOut[26] = fifoOut[45][14][w-1];
              unloadMuxOut[27] = fifoOut[46][14][w-1];
              unloadMuxOut[28] = fifoOut[47][14][w-1];
              unloadMuxOut[29] = fifoOut[48][14][w-1];
              unloadMuxOut[30] = fifoOut[49][14][w-1];
              unloadMuxOut[31] = fifoOut[50][14][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[51][15][w-1];
              unloadMuxOut[1] = fifoOut[26][14][w-1];
              unloadMuxOut[2] = fifoOut[27][14][w-1];
              unloadMuxOut[3] = fifoOut[28][14][w-1];
              unloadMuxOut[4] = fifoOut[29][14][w-1];
              unloadMuxOut[5] = fifoOut[30][14][w-1];
              unloadMuxOut[6] = fifoOut[31][14][w-1];
              unloadMuxOut[7] = fifoOut[32][14][w-1];
              unloadMuxOut[8] = fifoOut[33][14][w-1];
              unloadMuxOut[9] = fifoOut[34][14][w-1];
              unloadMuxOut[10] = fifoOut[35][14][w-1];
              unloadMuxOut[11] = fifoOut[36][14][w-1];
              unloadMuxOut[12] = fifoOut[37][14][w-1];
              unloadMuxOut[13] = fifoOut[38][14][w-1];
              unloadMuxOut[14] = fifoOut[39][14][w-1];
              unloadMuxOut[15] = fifoOut[40][14][w-1];
              unloadMuxOut[16] = fifoOut[41][14][w-1];
              unloadMuxOut[17] = fifoOut[42][14][w-1];
              unloadMuxOut[18] = fifoOut[43][14][w-1];
              unloadMuxOut[19] = fifoOut[44][14][w-1];
              unloadMuxOut[20] = fifoOut[45][14][w-1];
              unloadMuxOut[21] = fifoOut[46][14][w-1];
              unloadMuxOut[22] = fifoOut[47][14][w-1];
              unloadMuxOut[23] = fifoOut[48][14][w-1];
              unloadMuxOut[24] = fifoOut[49][14][w-1];
              unloadMuxOut[25] = fifoOut[50][14][w-1];
              unloadMuxOut[26] = fifoOut[51][14][w-1];
              unloadMuxOut[27] = fifoOut[26][13][w-1];
              unloadMuxOut[28] = fifoOut[27][13][w-1];
              unloadMuxOut[29] = fifoOut[28][13][w-1];
              unloadMuxOut[30] = fifoOut[29][13][w-1];
              unloadMuxOut[31] = fifoOut[30][13][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[31][14][w-1];
              unloadMuxOut[1] = fifoOut[32][14][w-1];
              unloadMuxOut[2] = fifoOut[33][14][w-1];
              unloadMuxOut[3] = fifoOut[34][14][w-1];
              unloadMuxOut[4] = fifoOut[35][14][w-1];
              unloadMuxOut[5] = fifoOut[36][14][w-1];
              unloadMuxOut[6] = fifoOut[37][14][w-1];
              unloadMuxOut[7] = fifoOut[38][14][w-1];
              unloadMuxOut[8] = fifoOut[39][14][w-1];
              unloadMuxOut[9] = fifoOut[40][14][w-1];
              unloadMuxOut[10] = fifoOut[41][14][w-1];
              unloadMuxOut[11] = fifoOut[42][14][w-1];
              unloadMuxOut[12] = fifoOut[43][14][w-1];
              unloadMuxOut[13] = fifoOut[44][14][w-1];
              unloadMuxOut[14] = fifoOut[45][14][w-1];
              unloadMuxOut[15] = fifoOut[46][14][w-1];
              unloadMuxOut[16] = fifoOut[47][14][w-1];
              unloadMuxOut[17] = fifoOut[48][14][w-1];
              unloadMuxOut[18] = fifoOut[49][14][w-1];
              unloadMuxOut[19] = fifoOut[50][14][w-1];
              unloadMuxOut[20] = fifoOut[51][14][w-1];
              unloadMuxOut[21] = fifoOut[26][13][w-1];
              unloadMuxOut[22] = fifoOut[27][13][w-1];
              unloadMuxOut[23] = fifoOut[28][13][w-1];
              unloadMuxOut[24] = fifoOut[29][13][w-1];
              unloadMuxOut[25] = fifoOut[30][13][w-1];
              unloadMuxOut[26] = fifoOut[31][13][w-1];
              unloadMuxOut[27] = fifoOut[32][13][w-1];
              unloadMuxOut[28] = fifoOut[33][13][w-1];
              unloadMuxOut[29] = fifoOut[34][13][w-1];
              unloadMuxOut[30] = fifoOut[35][13][w-1];
              unloadMuxOut[31] = fifoOut[36][13][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[37][14][w-1];
              unloadMuxOut[1] = fifoOut[38][14][w-1];
              unloadMuxOut[2] = fifoOut[39][14][w-1];
              unloadMuxOut[3] = fifoOut[40][14][w-1];
              unloadMuxOut[4] = fifoOut[41][14][w-1];
              unloadMuxOut[5] = fifoOut[42][14][w-1];
              unloadMuxOut[6] = fifoOut[43][14][w-1];
              unloadMuxOut[7] = fifoOut[44][14][w-1];
              unloadMuxOut[8] = fifoOut[45][14][w-1];
              unloadMuxOut[9] = fifoOut[46][14][w-1];
              unloadMuxOut[10] = fifoOut[47][14][w-1];
              unloadMuxOut[11] = fifoOut[48][14][w-1];
              unloadMuxOut[12] = fifoOut[49][14][w-1];
              unloadMuxOut[13] = fifoOut[50][14][w-1];
              unloadMuxOut[14] = fifoOut[51][14][w-1];
              unloadMuxOut[15] = fifoOut[26][13][w-1];
              unloadMuxOut[16] = fifoOut[27][13][w-1];
              unloadMuxOut[17] = fifoOut[28][13][w-1];
              unloadMuxOut[18] = fifoOut[29][13][w-1];
              unloadMuxOut[19] = fifoOut[30][13][w-1];
              unloadMuxOut[20] = fifoOut[31][13][w-1];
              unloadMuxOut[21] = fifoOut[32][13][w-1];
              unloadMuxOut[22] = fifoOut[33][13][w-1];
              unloadMuxOut[23] = fifoOut[34][13][w-1];
              unloadMuxOut[24] = fifoOut[35][13][w-1];
              unloadMuxOut[25] = fifoOut[36][13][w-1];
              unloadMuxOut[26] = fifoOut[37][13][w-1];
              unloadMuxOut[27] = fifoOut[38][13][w-1];
              unloadMuxOut[28] = fifoOut[39][13][w-1];
              unloadMuxOut[29] = fifoOut[40][13][w-1];
              unloadMuxOut[30] = fifoOut[41][13][w-1];
              unloadMuxOut[31] = fifoOut[42][13][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[23][9][w-1];
              unloadMuxOut[1] = fifoOut[24][9][w-1];
              unloadMuxOut[2] = fifoOut[25][9][w-1];
              unloadMuxOut[3] = fifoOut[0][8][w-1];
              unloadMuxOut[4] = fifoOut[1][8][w-1];
              unloadMuxOut[5] = fifoOut[2][8][w-1];
              unloadMuxOut[6] = fifoOut[3][8][w-1];
              unloadMuxOut[7] = fifoOut[4][8][w-1];
              unloadMuxOut[8] = fifoOut[5][8][w-1];
              unloadMuxOut[9] = fifoOut[6][8][w-1];
              unloadMuxOut[10] = fifoOut[7][8][w-1];
              unloadMuxOut[11] = fifoOut[8][8][w-1];
              unloadMuxOut[12] = fifoOut[9][8][w-1];
              unloadMuxOut[13] = fifoOut[10][8][w-1];
              unloadMuxOut[14] = fifoOut[11][8][w-1];
              unloadMuxOut[15] = fifoOut[12][8][w-1];
              unloadMuxOut[16] = fifoOut[13][8][w-1];
              unloadMuxOut[17] = fifoOut[14][8][w-1];
              unloadMuxOut[18] = fifoOut[15][8][w-1];
              unloadMuxOut[19] = fifoOut[16][8][w-1];
              unloadMuxOut[20] = fifoOut[17][8][w-1];
              unloadMuxOut[21] = fifoOut[18][8][w-1];
              unloadMuxOut[22] = fifoOut[19][8][w-1];
              unloadMuxOut[23] = fifoOut[20][8][w-1];
              unloadMuxOut[24] = fifoOut[21][8][w-1];
              unloadMuxOut[25] = fifoOut[22][8][w-1];
              unloadMuxOut[26] = fifoOut[23][8][w-1];
              unloadMuxOut[27] = fifoOut[24][8][w-1];
              unloadMuxOut[28] = fifoOut[25][8][w-1];
              unloadMuxOut[29] = fifoOut[0][7][w-1];
              unloadMuxOut[30] = fifoOut[1][7][w-1];
              unloadMuxOut[31] = fifoOut[2][7][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[3][8][w-1];
              unloadMuxOut[1] = fifoOut[4][8][w-1];
              unloadMuxOut[2] = fifoOut[5][8][w-1];
              unloadMuxOut[3] = fifoOut[6][8][w-1];
              unloadMuxOut[4] = fifoOut[7][8][w-1];
              unloadMuxOut[5] = fifoOut[8][8][w-1];
              unloadMuxOut[6] = fifoOut[9][8][w-1];
              unloadMuxOut[7] = fifoOut[10][8][w-1];
              unloadMuxOut[8] = fifoOut[11][8][w-1];
              unloadMuxOut[9] = fifoOut[12][8][w-1];
              unloadMuxOut[10] = fifoOut[13][8][w-1];
              unloadMuxOut[11] = fifoOut[14][8][w-1];
              unloadMuxOut[12] = fifoOut[15][8][w-1];
              unloadMuxOut[13] = fifoOut[16][8][w-1];
              unloadMuxOut[14] = fifoOut[17][8][w-1];
              unloadMuxOut[15] = fifoOut[18][8][w-1];
              unloadMuxOut[16] = fifoOut[19][8][w-1];
              unloadMuxOut[17] = fifoOut[20][8][w-1];
              unloadMuxOut[18] = fifoOut[21][8][w-1];
              unloadMuxOut[19] = fifoOut[22][8][w-1];
              unloadMuxOut[20] = fifoOut[23][8][w-1];
              unloadMuxOut[21] = fifoOut[24][8][w-1];
              unloadMuxOut[22] = fifoOut[25][8][w-1];
              unloadMuxOut[23] = fifoOut[0][7][w-1];
              unloadMuxOut[24] = fifoOut[1][7][w-1];
              unloadMuxOut[25] = fifoOut[2][7][w-1];
              unloadMuxOut[26] = fifoOut[3][7][w-1];
              unloadMuxOut[27] = fifoOut[4][7][w-1];
              unloadMuxOut[28] = fifoOut[5][7][w-1];
              unloadMuxOut[29] = fifoOut[6][7][w-1];
              unloadMuxOut[30] = fifoOut[7][7][w-1];
              unloadMuxOut[31] = fifoOut[8][7][w-1];
       end
       16: begin
              unloadMuxOut[0] = fifoOut[9][8][w-1];
              unloadMuxOut[1] = fifoOut[10][8][w-1];
              unloadMuxOut[2] = fifoOut[11][8][w-1];
              unloadMuxOut[3] = fifoOut[12][8][w-1];
              unloadMuxOut[4] = fifoOut[13][8][w-1];
              unloadMuxOut[5] = fifoOut[14][8][w-1];
              unloadMuxOut[6] = fifoOut[15][8][w-1];
              unloadMuxOut[7] = fifoOut[16][8][w-1];
              unloadMuxOut[8] = fifoOut[17][8][w-1];
              unloadMuxOut[9] = fifoOut[18][8][w-1];
              unloadMuxOut[10] = fifoOut[19][8][w-1];
              unloadMuxOut[11] = fifoOut[20][8][w-1];
              unloadMuxOut[12] = fifoOut[21][8][w-1];
              unloadMuxOut[13] = fifoOut[22][8][w-1];
              unloadMuxOut[14] = fifoOut[23][8][w-1];
              unloadMuxOut[15] = fifoOut[24][8][w-1];
              unloadMuxOut[16] = fifoOut[25][8][w-1];
              unloadMuxOut[17] = fifoOut[0][7][w-1];
              unloadMuxOut[18] = fifoOut[1][7][w-1];
              unloadMuxOut[19] = fifoOut[2][7][w-1];
              unloadMuxOut[20] = fifoOut[3][7][w-1];
              unloadMuxOut[21] = fifoOut[4][7][w-1];
              unloadMuxOut[22] = fifoOut[5][7][w-1];
              unloadMuxOut[23] = fifoOut[6][7][w-1];
              unloadMuxOut[24] = fifoOut[7][7][w-1];
              unloadMuxOut[25] = fifoOut[8][7][w-1];
              unloadMuxOut[26] = fifoOut[9][7][w-1];
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0; 
             end
       end
    endcase //unload case end
    case(iteration_0_indicator)
       0: begin
         case(rd_address_case)
         0: begin
              muxOutConnector[0] = fifoOut[10][8];
              muxOutConnector[1] = fifoOut[11][8];
              muxOutConnector[2] = fifoOut[12][8];
              muxOutConnector[3] = fifoOut[13][8];
              muxOutConnector[4] = fifoOut[14][8];
              muxOutConnector[5] = fifoOut[15][8];
              muxOutConnector[6] = fifoOut[16][8];
              muxOutConnector[7] = fifoOut[17][8];
              muxOutConnector[8] = fifoOut[18][8];
              muxOutConnector[9] = fifoOut[19][8];
              muxOutConnector[10] = fifoOut[20][8];
              muxOutConnector[11] = fifoOut[21][8];
              muxOutConnector[12] = fifoOut[22][8];
              muxOutConnector[13] = fifoOut[23][8];
              muxOutConnector[14] = fifoOut[24][8];
              muxOutConnector[15] = fifoOut[25][8];
              muxOutConnector[16] = fifoOut[0][7];
              muxOutConnector[17] = fifoOut[1][7];
              muxOutConnector[18] = fifoOut[2][7];
              muxOutConnector[19] = fifoOut[3][7];
              muxOutConnector[20] = fifoOut[4][7];
              muxOutConnector[21] = fifoOut[5][7];
              muxOutConnector[22] = fifoOut[6][7];
              muxOutConnector[23] = fifoOut[7][7];
              muxOutConnector[24] = fifoOut[8][7];
              muxOutConnector[25] = fifoOut[9][7];
              muxOutConnector[26] = fifoOut[41][1];
              muxOutConnector[27] = fifoOut[42][1];
              muxOutConnector[28] = fifoOut[43][1];
              muxOutConnector[29] = fifoOut[44][1];
              muxOutConnector[30] = fifoOut[45][1];
              muxOutConnector[31] = fifoOut[0][12];
              muxOutConnector[32] = fifoOut[1][12];
              muxOutConnector[33] = fifoOut[2][12];
              muxOutConnector[34] = fifoOut[3][12];
              muxOutConnector[35] = fifoOut[4][12];
              muxOutConnector[36] = fifoOut[5][12];
              muxOutConnector[37] = fifoOut[6][12];
              muxOutConnector[38] = fifoOut[7][12];
              muxOutConnector[39] = fifoOut[8][12];
              muxOutConnector[40] = fifoOut[9][12];
              muxOutConnector[41] = fifoOut[10][12];
              muxOutConnector[42] = fifoOut[11][12];
              muxOutConnector[43] = fifoOut[12][12];
              muxOutConnector[44] = fifoOut[13][12];
              muxOutConnector[45] = fifoOut[14][12];
              muxOutConnector[46] = fifoOut[15][12];
              muxOutConnector[47] = fifoOut[16][12];
              muxOutConnector[48] = fifoOut[17][12];
              muxOutConnector[49] = fifoOut[18][12];
              muxOutConnector[50] = fifoOut[19][12];
              muxOutConnector[51] = fifoOut[20][12];
         end
         1: begin
              muxOutConnector[0] = fifoOut[10][8];
              muxOutConnector[1] = fifoOut[11][8];
              muxOutConnector[2] = fifoOut[12][8];
              muxOutConnector[3] = fifoOut[13][8];
              muxOutConnector[4] = fifoOut[14][8];
              muxOutConnector[5] = fifoOut[15][8];
              muxOutConnector[6] = fifoOut[16][8];
              muxOutConnector[7] = fifoOut[17][8];
              muxOutConnector[8] = fifoOut[18][8];
              muxOutConnector[9] = fifoOut[19][8];
              muxOutConnector[10] = fifoOut[20][8];
              muxOutConnector[11] = fifoOut[21][8];
              muxOutConnector[12] = fifoOut[22][8];
              muxOutConnector[13] = fifoOut[23][8];
              muxOutConnector[14] = fifoOut[24][8];
              muxOutConnector[15] = fifoOut[25][8];
              muxOutConnector[16] = fifoOut[0][7];
              muxOutConnector[17] = fifoOut[1][7];
              muxOutConnector[18] = fifoOut[2][7];
              muxOutConnector[19] = fifoOut[3][7];
              muxOutConnector[20] = fifoOut[4][7];
              muxOutConnector[21] = fifoOut[5][7];
              muxOutConnector[22] = fifoOut[6][7];
              muxOutConnector[23] = fifoOut[7][7];
              muxOutConnector[24] = fifoOut[8][7];
              muxOutConnector[25] = fifoOut[9][7];
              muxOutConnector[26] = fifoOut[21][13];
              muxOutConnector[27] = fifoOut[22][13];
              muxOutConnector[28] = fifoOut[23][13];
              muxOutConnector[29] = fifoOut[24][13];
              muxOutConnector[30] = fifoOut[25][13];
              muxOutConnector[31] = fifoOut[0][12];
              muxOutConnector[32] = fifoOut[1][12];
              muxOutConnector[33] = fifoOut[2][12];
              muxOutConnector[34] = fifoOut[3][12];
              muxOutConnector[35] = fifoOut[4][12];
              muxOutConnector[36] = fifoOut[5][12];
              muxOutConnector[37] = fifoOut[6][12];
              muxOutConnector[38] = fifoOut[7][12];
              muxOutConnector[39] = fifoOut[8][12];
              muxOutConnector[40] = fifoOut[9][12];
              muxOutConnector[41] = fifoOut[10][12];
              muxOutConnector[42] = fifoOut[11][12];
              muxOutConnector[43] = fifoOut[12][12];
              muxOutConnector[44] = fifoOut[13][12];
              muxOutConnector[45] = fifoOut[14][12];
              muxOutConnector[46] = fifoOut[15][12];
              muxOutConnector[47] = fifoOut[16][12];
              muxOutConnector[48] = fifoOut[17][12];
              muxOutConnector[49] = fifoOut[18][12];
              muxOutConnector[50] = fifoOut[19][12];
              muxOutConnector[51] = fifoOut[20][12];
         end
         2: begin
              muxOutConnector[0] = fifoOut[10][8];
              muxOutConnector[1] = fifoOut[11][8];
              muxOutConnector[2] = fifoOut[12][8];
              muxOutConnector[3] = fifoOut[13][8];
              muxOutConnector[4] = fifoOut[14][8];
              muxOutConnector[5] = fifoOut[15][8];
              muxOutConnector[6] = fifoOut[16][8];
              muxOutConnector[7] = fifoOut[17][8];
              muxOutConnector[8] = fifoOut[18][8];
              muxOutConnector[9] = fifoOut[19][8];
              muxOutConnector[10] = fifoOut[20][8];
              muxOutConnector[11] = fifoOut[21][8];
              muxOutConnector[12] = fifoOut[22][8];
              muxOutConnector[13] = fifoOut[23][8];
              muxOutConnector[14] = fifoOut[24][8];
              muxOutConnector[15] = fifoOut[25][8];
              muxOutConnector[16] = fifoOut[0][7];
              muxOutConnector[17] = fifoOut[1][7];
              muxOutConnector[18] = fifoOut[2][7];
              muxOutConnector[19] = fifoOut[3][7];
              muxOutConnector[20] = fifoOut[4][7];
              muxOutConnector[21] = fifoOut[5][7];
              muxOutConnector[22] = fifoOut[6][7];
              muxOutConnector[23] = fifoOut[7][7];
              muxOutConnector[24] = fifoOut[8][7];
              muxOutConnector[25] = fifoOut[9][7];
              muxOutConnector[26] = fifoOut[21][13];
              muxOutConnector[27] = fifoOut[22][13];
              muxOutConnector[28] = fifoOut[23][13];
              muxOutConnector[29] = fifoOut[24][13];
              muxOutConnector[30] = fifoOut[25][13];
              muxOutConnector[31] = fifoOut[0][12];
              muxOutConnector[32] = fifoOut[1][12];
              muxOutConnector[33] = fifoOut[2][12];
              muxOutConnector[34] = fifoOut[3][12];
              muxOutConnector[35] = fifoOut[4][12];
              muxOutConnector[36] = fifoOut[5][12];
              muxOutConnector[37] = fifoOut[6][12];
              muxOutConnector[38] = fifoOut[7][12];
              muxOutConnector[39] = fifoOut[8][12];
              muxOutConnector[40] = fifoOut[9][12];
              muxOutConnector[41] = fifoOut[10][12];
              muxOutConnector[42] = fifoOut[11][12];
              muxOutConnector[43] = fifoOut[12][12];
              muxOutConnector[44] = fifoOut[13][12];
              muxOutConnector[45] = fifoOut[14][12];
              muxOutConnector[46] = fifoOut[15][12];
              muxOutConnector[47] = fifoOut[16][12];
              muxOutConnector[48] = fifoOut[17][12];
              muxOutConnector[49] = fifoOut[18][12];
              muxOutConnector[50] = fifoOut[19][12];
              muxOutConnector[51] = fifoOut[20][12];
         end
         3: begin
              muxOutConnector[0] = fifoOut[10][8];
              muxOutConnector[1] = fifoOut[11][8];
              muxOutConnector[2] = fifoOut[12][8];
              muxOutConnector[3] = fifoOut[13][8];
              muxOutConnector[4] = fifoOut[14][8];
              muxOutConnector[5] = fifoOut[15][8];
              muxOutConnector[6] = fifoOut[16][8];
              muxOutConnector[7] = fifoOut[17][8];
              muxOutConnector[8] = fifoOut[18][8];
              muxOutConnector[9] = fifoOut[19][8];
              muxOutConnector[10] = fifoOut[20][8];
              muxOutConnector[11] = fifoOut[21][8];
              muxOutConnector[12] = fifoOut[22][8];
              muxOutConnector[13] = fifoOut[26][15];
              muxOutConnector[14] = fifoOut[27][15];
              muxOutConnector[15] = fifoOut[28][15];
              muxOutConnector[16] = fifoOut[29][15];
              muxOutConnector[17] = fifoOut[30][15];
              muxOutConnector[18] = fifoOut[31][15];
              muxOutConnector[19] = fifoOut[32][15];
              muxOutConnector[20] = fifoOut[33][15];
              muxOutConnector[21] = fifoOut[34][15];
              muxOutConnector[22] = fifoOut[35][15];
              muxOutConnector[23] = fifoOut[36][15];
              muxOutConnector[24] = fifoOut[37][15];
              muxOutConnector[25] = fifoOut[38][15];
              muxOutConnector[26] = fifoOut[21][13];
              muxOutConnector[27] = fifoOut[22][13];
              muxOutConnector[28] = fifoOut[23][13];
              muxOutConnector[29] = fifoOut[24][13];
              muxOutConnector[30] = fifoOut[25][13];
              muxOutConnector[31] = fifoOut[0][12];
              muxOutConnector[32] = fifoOut[1][12];
              muxOutConnector[33] = fifoOut[2][12];
              muxOutConnector[34] = fifoOut[3][12];
              muxOutConnector[35] = fifoOut[4][12];
              muxOutConnector[36] = fifoOut[5][12];
              muxOutConnector[37] = fifoOut[6][12];
              muxOutConnector[38] = fifoOut[7][12];
              muxOutConnector[39] = fifoOut[8][12];
              muxOutConnector[40] = fifoOut[9][12];
              muxOutConnector[41] = fifoOut[10][12];
              muxOutConnector[42] = fifoOut[11][12];
              muxOutConnector[43] = fifoOut[12][12];
              muxOutConnector[44] = fifoOut[13][12];
              muxOutConnector[45] = fifoOut[14][12];
              muxOutConnector[46] = fifoOut[15][12];
              muxOutConnector[47] = fifoOut[16][12];
              muxOutConnector[48] = fifoOut[17][12];
              muxOutConnector[49] = fifoOut[18][12];
              muxOutConnector[50] = fifoOut[19][12];
              muxOutConnector[51] = fifoOut[20][12];
         end
         4: begin
              muxOutConnector[0] = fifoOut[39][16];
              muxOutConnector[1] = fifoOut[40][16];
              muxOutConnector[2] = fifoOut[41][16];
              muxOutConnector[3] = fifoOut[42][16];
              muxOutConnector[4] = fifoOut[43][16];
              muxOutConnector[5] = fifoOut[44][16];
              muxOutConnector[6] = fifoOut[45][16];
              muxOutConnector[7] = fifoOut[46][16];
              muxOutConnector[8] = fifoOut[47][16];
              muxOutConnector[9] = fifoOut[48][16];
              muxOutConnector[10] = fifoOut[49][16];
              muxOutConnector[11] = fifoOut[50][16];
              muxOutConnector[12] = fifoOut[51][16];
              muxOutConnector[13] = fifoOut[26][15];
              muxOutConnector[14] = fifoOut[27][15];
              muxOutConnector[15] = fifoOut[28][15];
              muxOutConnector[16] = fifoOut[29][15];
              muxOutConnector[17] = fifoOut[30][15];
              muxOutConnector[18] = fifoOut[31][15];
              muxOutConnector[19] = fifoOut[32][15];
              muxOutConnector[20] = fifoOut[33][15];
              muxOutConnector[21] = fifoOut[34][15];
              muxOutConnector[22] = fifoOut[35][15];
              muxOutConnector[23] = fifoOut[36][15];
              muxOutConnector[24] = fifoOut[37][15];
              muxOutConnector[25] = fifoOut[38][15];
              muxOutConnector[26] = fifoOut[21][13];
              muxOutConnector[27] = fifoOut[22][13];
              muxOutConnector[28] = fifoOut[23][13];
              muxOutConnector[29] = fifoOut[24][13];
              muxOutConnector[30] = fifoOut[25][13];
              muxOutConnector[31] = fifoOut[0][12];
              muxOutConnector[32] = fifoOut[1][12];
              muxOutConnector[33] = fifoOut[2][12];
              muxOutConnector[34] = fifoOut[3][12];
              muxOutConnector[35] = fifoOut[4][12];
              muxOutConnector[36] = fifoOut[5][12];
              muxOutConnector[37] = fifoOut[6][12];
              muxOutConnector[38] = fifoOut[7][12];
              muxOutConnector[39] = fifoOut[8][12];
              muxOutConnector[40] = fifoOut[9][12];
              muxOutConnector[41] = fifoOut[10][12];
              muxOutConnector[42] = fifoOut[11][12];
              muxOutConnector[43] = fifoOut[12][12];
              muxOutConnector[44] = fifoOut[13][12];
              muxOutConnector[45] = fifoOut[14][12];
              muxOutConnector[46] = fifoOut[15][12];
              muxOutConnector[47] = fifoOut[16][12];
              muxOutConnector[48] = fifoOut[17][12];
              muxOutConnector[49] = fifoOut[18][12];
              muxOutConnector[50] = fifoOut[19][12];
              muxOutConnector[51] = fifoOut[20][12];
         end
         5: begin
              muxOutConnector[0] = fifoOut[39][16];
              muxOutConnector[1] = fifoOut[40][16];
              muxOutConnector[2] = fifoOut[41][16];
              muxOutConnector[3] = fifoOut[42][16];
              muxOutConnector[4] = fifoOut[43][16];
              muxOutConnector[5] = fifoOut[44][16];
              muxOutConnector[6] = fifoOut[45][16];
              muxOutConnector[7] = fifoOut[46][16];
              muxOutConnector[8] = fifoOut[47][16];
              muxOutConnector[9] = fifoOut[48][16];
              muxOutConnector[10] = fifoOut[49][16];
              muxOutConnector[11] = fifoOut[50][16];
              muxOutConnector[12] = fifoOut[51][16];
              muxOutConnector[13] = fifoOut[26][15];
              muxOutConnector[14] = fifoOut[27][15];
              muxOutConnector[15] = fifoOut[28][15];
              muxOutConnector[16] = fifoOut[29][15];
              muxOutConnector[17] = fifoOut[30][15];
              muxOutConnector[18] = fifoOut[31][15];
              muxOutConnector[19] = fifoOut[32][15];
              muxOutConnector[20] = fifoOut[33][15];
              muxOutConnector[21] = fifoOut[34][15];
              muxOutConnector[22] = fifoOut[35][15];
              muxOutConnector[23] = fifoOut[36][15];
              muxOutConnector[24] = fifoOut[37][15];
              muxOutConnector[25] = fifoOut[38][15];
              muxOutConnector[26] = fifoOut[21][13];
              muxOutConnector[27] = fifoOut[22][13];
              muxOutConnector[28] = fifoOut[23][13];
              muxOutConnector[29] = fifoOut[24][13];
              muxOutConnector[30] = fifoOut[25][13];
              muxOutConnector[31] = fifoOut[0][12];
              muxOutConnector[32] = fifoOut[1][12];
              muxOutConnector[33] = fifoOut[2][12];
              muxOutConnector[34] = fifoOut[3][12];
              muxOutConnector[35] = fifoOut[4][12];
              muxOutConnector[36] = fifoOut[5][12];
              muxOutConnector[37] = fifoOut[6][12];
              muxOutConnector[38] = fifoOut[7][12];
              muxOutConnector[39] = fifoOut[8][12];
              muxOutConnector[40] = fifoOut[9][12];
              muxOutConnector[41] = fifoOut[10][12];
              muxOutConnector[42] = fifoOut[11][12];
              muxOutConnector[43] = fifoOut[12][12];
              muxOutConnector[44] = fifoOut[13][12];
              muxOutConnector[45] = fifoOut[14][12];
              muxOutConnector[46] = fifoOut[15][12];
              muxOutConnector[47] = fifoOut[16][12];
              muxOutConnector[48] = fifoOut[17][12];
              muxOutConnector[49] = fifoOut[18][12];
              muxOutConnector[50] = fifoOut[19][12];
              muxOutConnector[51] = fifoOut[20][12];
         end
         6: begin
              muxOutConnector[0] = fifoOut[39][16];
              muxOutConnector[1] = fifoOut[40][16];
              muxOutConnector[2] = fifoOut[41][16];
              muxOutConnector[3] = fifoOut[42][16];
              muxOutConnector[4] = fifoOut[43][16];
              muxOutConnector[5] = fifoOut[44][16];
              muxOutConnector[6] = fifoOut[45][16];
              muxOutConnector[7] = fifoOut[46][16];
              muxOutConnector[8] = fifoOut[47][16];
              muxOutConnector[9] = fifoOut[48][16];
              muxOutConnector[10] = fifoOut[49][16];
              muxOutConnector[11] = fifoOut[50][16];
              muxOutConnector[12] = fifoOut[51][16];
              muxOutConnector[13] = fifoOut[26][15];
              muxOutConnector[14] = fifoOut[27][15];
              muxOutConnector[15] = fifoOut[28][15];
              muxOutConnector[16] = fifoOut[29][15];
              muxOutConnector[17] = fifoOut[30][15];
              muxOutConnector[18] = fifoOut[31][15];
              muxOutConnector[19] = fifoOut[32][15];
              muxOutConnector[20] = fifoOut[33][15];
              muxOutConnector[21] = fifoOut[34][15];
              muxOutConnector[22] = fifoOut[35][15];
              muxOutConnector[23] = fifoOut[36][15];
              muxOutConnector[24] = fifoOut[37][15];
              muxOutConnector[25] = fifoOut[38][15];
              muxOutConnector[26] = fifoOut[21][13];
              muxOutConnector[27] = fifoOut[22][13];
              muxOutConnector[28] = fifoOut[23][13];
              muxOutConnector[29] = fifoOut[24][13];
              muxOutConnector[30] = fifoOut[25][13];
              muxOutConnector[31] = fifoOut[0][12];
              muxOutConnector[32] = fifoOut[1][12];
              muxOutConnector[33] = fifoOut[2][12];
              muxOutConnector[34] = fifoOut[3][12];
              muxOutConnector[35] = fifoOut[4][12];
              muxOutConnector[36] = fifoOut[5][12];
              muxOutConnector[37] = fifoOut[6][12];
              muxOutConnector[38] = fifoOut[7][12];
              muxOutConnector[39] = fifoOut[8][12];
              muxOutConnector[40] = fifoOut[9][12];
              muxOutConnector[41] = fifoOut[10][12];
              muxOutConnector[42] = fifoOut[11][12];
              muxOutConnector[43] = fifoOut[12][12];
              muxOutConnector[44] = fifoOut[13][12];
              muxOutConnector[45] = fifoOut[14][12];
              muxOutConnector[46] = fifoOut[15][12];
              muxOutConnector[47] = fifoOut[16][12];
              muxOutConnector[48] = fifoOut[17][12];
              muxOutConnector[49] = fifoOut[18][12];
              muxOutConnector[50] = fifoOut[19][12];
              muxOutConnector[51] = fifoOut[20][12];
         end
         7: begin
              muxOutConnector[0] = fifoOut[39][16];
              muxOutConnector[1] = fifoOut[40][16];
              muxOutConnector[2] = fifoOut[41][16];
              muxOutConnector[3] = fifoOut[42][16];
              muxOutConnector[4] = fifoOut[43][16];
              muxOutConnector[5] = fifoOut[44][16];
              muxOutConnector[6] = fifoOut[45][16];
              muxOutConnector[7] = fifoOut[46][16];
              muxOutConnector[8] = fifoOut[47][16];
              muxOutConnector[9] = fifoOut[48][16];
              muxOutConnector[10] = fifoOut[49][16];
              muxOutConnector[11] = fifoOut[50][16];
              muxOutConnector[12] = fifoOut[51][16];
              muxOutConnector[13] = fifoOut[26][15];
              muxOutConnector[14] = fifoOut[27][15];
              muxOutConnector[15] = fifoOut[28][15];
              muxOutConnector[16] = fifoOut[29][15];
              muxOutConnector[17] = fifoOut[30][15];
              muxOutConnector[18] = fifoOut[31][15];
              muxOutConnector[19] = fifoOut[32][15];
              muxOutConnector[20] = fifoOut[33][15];
              muxOutConnector[21] = fifoOut[34][15];
              muxOutConnector[22] = fifoOut[35][15];
              muxOutConnector[23] = fifoOut[36][15];
              muxOutConnector[24] = fifoOut[37][15];
              muxOutConnector[25] = fifoOut[38][15];
              muxOutConnector[26] = fifoOut[21][13];
              muxOutConnector[27] = fifoOut[22][13];
              muxOutConnector[28] = fifoOut[23][13];
              muxOutConnector[29] = fifoOut[24][13];
              muxOutConnector[30] = fifoOut[25][13];
              muxOutConnector[31] = fifoOut[0][12];
              muxOutConnector[32] = fifoOut[1][12];
              muxOutConnector[33] = fifoOut[2][12];
              muxOutConnector[34] = fifoOut[3][12];
              muxOutConnector[35] = fifoOut[4][12];
              muxOutConnector[36] = fifoOut[5][12];
              muxOutConnector[37] = fifoOut[6][12];
              muxOutConnector[38] = fifoOut[7][12];
              muxOutConnector[39] = fifoOut[8][12];
              muxOutConnector[40] = fifoOut[9][12];
              muxOutConnector[41] = fifoOut[10][12];
              muxOutConnector[42] = fifoOut[11][12];
              muxOutConnector[43] = fifoOut[12][12];
              muxOutConnector[44] = fifoOut[13][12];
              muxOutConnector[45] = fifoOut[14][12];
              muxOutConnector[46] = fifoOut[15][12];
              muxOutConnector[47] = fifoOut[16][12];
              muxOutConnector[48] = fifoOut[17][12];
              muxOutConnector[49] = fifoOut[18][12];
              muxOutConnector[50] = fifoOut[19][12];
              muxOutConnector[51] = fifoOut[20][12];
         end
         8: begin
              muxOutConnector[0] = fifoOut[39][16];
              muxOutConnector[1] = fifoOut[40][16];
              muxOutConnector[2] = fifoOut[41][16];
              muxOutConnector[3] = fifoOut[42][16];
              muxOutConnector[4] = fifoOut[43][16];
              muxOutConnector[5] = fifoOut[44][16];
              muxOutConnector[6] = fifoOut[45][16];
              muxOutConnector[7] = fifoOut[46][16];
              muxOutConnector[8] = fifoOut[47][16];
              muxOutConnector[9] = fifoOut[48][16];
              muxOutConnector[10] = fifoOut[49][16];
              muxOutConnector[11] = fifoOut[50][16];
              muxOutConnector[12] = fifoOut[51][16];
              muxOutConnector[13] = fifoOut[26][15];
              muxOutConnector[14] = fifoOut[27][15];
              muxOutConnector[15] = fifoOut[28][15];
              muxOutConnector[16] = fifoOut[29][15];
              muxOutConnector[17] = fifoOut[30][15];
              muxOutConnector[18] = fifoOut[31][15];
              muxOutConnector[19] = fifoOut[32][15];
              muxOutConnector[20] = fifoOut[33][15];
              muxOutConnector[21] = fifoOut[34][15];
              muxOutConnector[22] = fifoOut[35][15];
              muxOutConnector[23] = fifoOut[36][15];
              muxOutConnector[24] = fifoOut[37][15];
              muxOutConnector[25] = fifoOut[38][15];
              muxOutConnector[26] = fifoOut[21][13];
              muxOutConnector[27] = fifoOut[22][13];
              muxOutConnector[28] = fifoOut[23][13];
              muxOutConnector[29] = fifoOut[24][13];
              muxOutConnector[30] = fifoOut[25][13];
              muxOutConnector[31] = fifoOut[0][12];
              muxOutConnector[32] = fifoOut[1][12];
              muxOutConnector[33] = fifoOut[2][12];
              muxOutConnector[34] = fifoOut[3][12];
              muxOutConnector[35] = fifoOut[4][12];
              muxOutConnector[36] = fifoOut[5][12];
              muxOutConnector[37] = fifoOut[6][12];
              muxOutConnector[38] = fifoOut[7][12];
              muxOutConnector[39] = fifoOut[8][12];
              muxOutConnector[40] = fifoOut[9][12];
              muxOutConnector[41] = fifoOut[10][12];
              muxOutConnector[42] = fifoOut[11][12];
              muxOutConnector[43] = fifoOut[12][12];
              muxOutConnector[44] = fifoOut[13][12];
              muxOutConnector[45] = fifoOut[14][12];
              muxOutConnector[46] = fifoOut[15][12];
              muxOutConnector[47] = fifoOut[16][12];
              muxOutConnector[48] = fifoOut[17][12];
              muxOutConnector[49] = fifoOut[18][12];
              muxOutConnector[50] = fifoOut[19][12];
              muxOutConnector[51] = fifoOut[20][12];
         end
         9: begin
              muxOutConnector[0] = fifoOut[39][16];
              muxOutConnector[1] = fifoOut[40][16];
              muxOutConnector[2] = fifoOut[41][16];
              muxOutConnector[3] = fifoOut[42][16];
              muxOutConnector[4] = fifoOut[43][16];
              muxOutConnector[5] = fifoOut[44][16];
              muxOutConnector[6] = fifoOut[45][16];
              muxOutConnector[7] = fifoOut[46][16];
              muxOutConnector[8] = fifoOut[47][16];
              muxOutConnector[9] = fifoOut[48][16];
              muxOutConnector[10] = fifoOut[49][16];
              muxOutConnector[11] = fifoOut[50][16];
              muxOutConnector[12] = fifoOut[51][16];
              muxOutConnector[13] = fifoOut[26][15];
              muxOutConnector[14] = fifoOut[27][15];
              muxOutConnector[15] = fifoOut[28][15];
              muxOutConnector[16] = fifoOut[29][15];
              muxOutConnector[17] = fifoOut[30][15];
              muxOutConnector[18] = fifoOut[31][15];
              muxOutConnector[19] = fifoOut[32][15];
              muxOutConnector[20] = fifoOut[33][15];
              muxOutConnector[21] = fifoOut[34][15];
              muxOutConnector[22] = fifoOut[35][15];
              muxOutConnector[23] = fifoOut[36][15];
              muxOutConnector[24] = fifoOut[37][15];
              muxOutConnector[25] = fifoOut[38][15];
              muxOutConnector[26] = fifoOut[21][13];
              muxOutConnector[27] = fifoOut[22][13];
              muxOutConnector[28] = fifoOut[23][13];
              muxOutConnector[29] = fifoOut[24][13];
              muxOutConnector[30] = fifoOut[25][13];
              muxOutConnector[31] = fifoOut[0][12];
              muxOutConnector[32] = fifoOut[1][12];
              muxOutConnector[33] = fifoOut[2][12];
              muxOutConnector[34] = fifoOut[3][12];
              muxOutConnector[35] = fifoOut[4][12];
              muxOutConnector[36] = fifoOut[5][12];
              muxOutConnector[37] = fifoOut[6][12];
              muxOutConnector[38] = fifoOut[7][12];
              muxOutConnector[39] = fifoOut[8][12];
              muxOutConnector[40] = fifoOut[9][12];
              muxOutConnector[41] = fifoOut[10][12];
              muxOutConnector[42] = fifoOut[11][12];
              muxOutConnector[43] = fifoOut[12][12];
              muxOutConnector[44] = fifoOut[13][12];
              muxOutConnector[45] = fifoOut[14][12];
              muxOutConnector[46] = fifoOut[15][12];
              muxOutConnector[47] = fifoOut[16][12];
              muxOutConnector[48] = fifoOut[17][12];
              muxOutConnector[49] = fifoOut[18][12];
              muxOutConnector[50] = fifoOut[19][12];
              muxOutConnector[51] = fifoOut[20][12];
         end
         10: begin
              muxOutConnector[0] = fifoOut[39][16];
              muxOutConnector[1] = fifoOut[40][16];
              muxOutConnector[2] = fifoOut[41][16];
              muxOutConnector[3] = fifoOut[42][16];
              muxOutConnector[4] = fifoOut[43][16];
              muxOutConnector[5] = fifoOut[44][16];
              muxOutConnector[6] = fifoOut[45][16];
              muxOutConnector[7] = fifoOut[46][16];
              muxOutConnector[8] = fifoOut[47][16];
              muxOutConnector[9] = fifoOut[48][16];
              muxOutConnector[10] = fifoOut[49][16];
              muxOutConnector[11] = fifoOut[50][16];
              muxOutConnector[12] = fifoOut[51][16];
              muxOutConnector[13] = fifoOut[26][15];
              muxOutConnector[14] = fifoOut[27][15];
              muxOutConnector[15] = fifoOut[28][15];
              muxOutConnector[16] = fifoOut[29][15];
              muxOutConnector[17] = fifoOut[30][15];
              muxOutConnector[18] = fifoOut[31][15];
              muxOutConnector[19] = fifoOut[32][15];
              muxOutConnector[20] = fifoOut[33][15];
              muxOutConnector[21] = fifoOut[34][15];
              muxOutConnector[22] = fifoOut[35][15];
              muxOutConnector[23] = fifoOut[36][15];
              muxOutConnector[24] = fifoOut[37][15];
              muxOutConnector[25] = fifoOut[38][15];
              muxOutConnector[26] = fifoOut[21][13];
              muxOutConnector[27] = fifoOut[22][13];
              muxOutConnector[28] = fifoOut[23][13];
              muxOutConnector[29] = fifoOut[24][13];
              muxOutConnector[30] = fifoOut[25][13];
              muxOutConnector[31] = fifoOut[0][12];
              muxOutConnector[32] = fifoOut[1][12];
              muxOutConnector[33] = fifoOut[2][12];
              muxOutConnector[34] = fifoOut[3][12];
              muxOutConnector[35] = fifoOut[4][12];
              muxOutConnector[36] = fifoOut[5][12];
              muxOutConnector[37] = fifoOut[6][12];
              muxOutConnector[38] = fifoOut[7][12];
              muxOutConnector[39] = fifoOut[8][12];
              muxOutConnector[40] = fifoOut[9][12];
              muxOutConnector[41] = fifoOut[10][12];
              muxOutConnector[42] = fifoOut[11][12];
              muxOutConnector[43] = fifoOut[12][12];
              muxOutConnector[44] = fifoOut[13][12];
              muxOutConnector[45] = fifoOut[14][12];
              muxOutConnector[46] = fifoOut[15][12];
              muxOutConnector[47] = fifoOut[16][12];
              muxOutConnector[48] = fifoOut[17][12];
              muxOutConnector[49] = fifoOut[18][12];
              muxOutConnector[50] = fifoOut[19][12];
              muxOutConnector[51] = fifoOut[20][12];
         end
         11: begin
              muxOutConnector[0] = fifoOut[39][16];
              muxOutConnector[1] = fifoOut[40][16];
              muxOutConnector[2] = fifoOut[41][16];
              muxOutConnector[3] = fifoOut[42][16];
              muxOutConnector[4] = fifoOut[43][16];
              muxOutConnector[5] = fifoOut[44][16];
              muxOutConnector[6] = fifoOut[45][16];
              muxOutConnector[7] = fifoOut[46][16];
              muxOutConnector[8] = fifoOut[47][16];
              muxOutConnector[9] = fifoOut[48][16];
              muxOutConnector[10] = fifoOut[49][16];
              muxOutConnector[11] = fifoOut[50][16];
              muxOutConnector[12] = fifoOut[51][16];
              muxOutConnector[13] = fifoOut[26][15];
              muxOutConnector[14] = fifoOut[27][15];
              muxOutConnector[15] = fifoOut[28][15];
              muxOutConnector[16] = fifoOut[29][15];
              muxOutConnector[17] = fifoOut[30][15];
              muxOutConnector[18] = fifoOut[31][15];
              muxOutConnector[19] = fifoOut[32][15];
              muxOutConnector[20] = fifoOut[33][15];
              muxOutConnector[21] = fifoOut[34][15];
              muxOutConnector[22] = fifoOut[35][15];
              muxOutConnector[23] = fifoOut[36][15];
              muxOutConnector[24] = fifoOut[37][15];
              muxOutConnector[25] = fifoOut[38][15];
              muxOutConnector[26] = fifoOut[21][13];
              muxOutConnector[27] = fifoOut[22][13];
              muxOutConnector[28] = fifoOut[23][13];
              muxOutConnector[29] = fifoOut[24][13];
              muxOutConnector[30] = fifoOut[25][13];
              muxOutConnector[31] = fifoOut[0][12];
              muxOutConnector[32] = fifoOut[1][12];
              muxOutConnector[33] = fifoOut[2][12];
              muxOutConnector[34] = fifoOut[3][12];
              muxOutConnector[35] = fifoOut[4][12];
              muxOutConnector[36] = fifoOut[5][12];
              muxOutConnector[37] = fifoOut[6][12];
              muxOutConnector[38] = fifoOut[7][12];
              muxOutConnector[39] = fifoOut[8][12];
              muxOutConnector[40] = fifoOut[9][12];
              muxOutConnector[41] = fifoOut[10][12];
              muxOutConnector[42] = fifoOut[11][12];
              muxOutConnector[43] = fifoOut[12][12];
              muxOutConnector[44] = fifoOut[13][12];
              muxOutConnector[45] = fifoOut[14][12];
              muxOutConnector[46] = fifoOut[15][12];
              muxOutConnector[47] = fifoOut[16][12];
              muxOutConnector[48] = fifoOut[17][12];
              muxOutConnector[49] = fifoOut[18][12];
              muxOutConnector[50] = fifoOut[19][12];
              muxOutConnector[51] = fifoOut[20][12];
         end
         12: begin
              muxOutConnector[0] = fifoOut[39][16];
              muxOutConnector[1] = fifoOut[40][16];
              muxOutConnector[2] = fifoOut[41][16];
              muxOutConnector[3] = fifoOut[42][16];
              muxOutConnector[4] = fifoOut[43][16];
              muxOutConnector[5] = fifoOut[44][16];
              muxOutConnector[6] = fifoOut[45][16];
              muxOutConnector[7] = fifoOut[46][16];
              muxOutConnector[8] = fifoOut[47][16];
              muxOutConnector[9] = fifoOut[48][16];
              muxOutConnector[10] = fifoOut[49][16];
              muxOutConnector[11] = fifoOut[50][16];
              muxOutConnector[12] = fifoOut[51][16];
              muxOutConnector[13] = fifoOut[26][15];
              muxOutConnector[14] = fifoOut[27][15];
              muxOutConnector[15] = fifoOut[28][15];
              muxOutConnector[16] = fifoOut[29][15];
              muxOutConnector[17] = fifoOut[30][15];
              muxOutConnector[18] = fifoOut[31][15];
              muxOutConnector[19] = fifoOut[32][15];
              muxOutConnector[20] = fifoOut[33][15];
              muxOutConnector[21] = fifoOut[34][15];
              muxOutConnector[22] = fifoOut[35][15];
              muxOutConnector[23] = fifoOut[36][15];
              muxOutConnector[24] = fifoOut[37][15];
              muxOutConnector[25] = fifoOut[38][15];
              muxOutConnector[26] = fifoOut[21][13];
              muxOutConnector[27] = fifoOut[22][13];
              muxOutConnector[28] = fifoOut[23][13];
              muxOutConnector[29] = fifoOut[24][13];
              muxOutConnector[30] = fifoOut[25][13];
              muxOutConnector[31] = fifoOut[0][12];
              muxOutConnector[32] = fifoOut[1][12];
              muxOutConnector[33] = fifoOut[2][12];
              muxOutConnector[34] = fifoOut[3][12];
              muxOutConnector[35] = fifoOut[4][12];
              muxOutConnector[36] = fifoOut[5][12];
              muxOutConnector[37] = fifoOut[6][12];
              muxOutConnector[38] = fifoOut[7][12];
              muxOutConnector[39] = fifoOut[8][12];
              muxOutConnector[40] = fifoOut[9][12];
              muxOutConnector[41] = fifoOut[10][12];
              muxOutConnector[42] = fifoOut[11][12];
              muxOutConnector[43] = fifoOut[12][12];
              muxOutConnector[44] = fifoOut[13][12];
              muxOutConnector[45] = fifoOut[14][12];
              muxOutConnector[46] = fifoOut[15][12];
              muxOutConnector[47] = fifoOut[16][12];
              muxOutConnector[48] = fifoOut[46][3];
              muxOutConnector[49] = fifoOut[47][3];
              muxOutConnector[50] = fifoOut[48][3];
              muxOutConnector[51] = fifoOut[49][3];
         end
         13: begin
              muxOutConnector[0] = fifoOut[39][16];
              muxOutConnector[1] = fifoOut[40][16];
              muxOutConnector[2] = fifoOut[41][16];
              muxOutConnector[3] = fifoOut[42][16];
              muxOutConnector[4] = fifoOut[43][16];
              muxOutConnector[5] = fifoOut[44][16];
              muxOutConnector[6] = fifoOut[45][16];
              muxOutConnector[7] = fifoOut[46][16];
              muxOutConnector[8] = fifoOut[47][16];
              muxOutConnector[9] = fifoOut[48][16];
              muxOutConnector[10] = fifoOut[49][16];
              muxOutConnector[11] = fifoOut[50][16];
              muxOutConnector[12] = fifoOut[51][16];
              muxOutConnector[13] = fifoOut[26][15];
              muxOutConnector[14] = fifoOut[27][15];
              muxOutConnector[15] = fifoOut[28][15];
              muxOutConnector[16] = fifoOut[29][15];
              muxOutConnector[17] = fifoOut[30][15];
              muxOutConnector[18] = fifoOut[31][15];
              muxOutConnector[19] = fifoOut[32][15];
              muxOutConnector[20] = fifoOut[33][15];
              muxOutConnector[21] = fifoOut[34][15];
              muxOutConnector[22] = fifoOut[35][15];
              muxOutConnector[23] = fifoOut[36][15];
              muxOutConnector[24] = fifoOut[37][15];
              muxOutConnector[25] = fifoOut[38][15];
              muxOutConnector[26] = fifoOut[50][4];
              muxOutConnector[27] = fifoOut[51][4];
              muxOutConnector[28] = fifoOut[26][3];
              muxOutConnector[29] = fifoOut[27][3];
              muxOutConnector[30] = fifoOut[28][3];
              muxOutConnector[31] = fifoOut[29][3];
              muxOutConnector[32] = fifoOut[30][3];
              muxOutConnector[33] = fifoOut[31][3];
              muxOutConnector[34] = fifoOut[32][3];
              muxOutConnector[35] = fifoOut[33][3];
              muxOutConnector[36] = fifoOut[34][3];
              muxOutConnector[37] = fifoOut[35][3];
              muxOutConnector[38] = fifoOut[36][3];
              muxOutConnector[39] = fifoOut[37][3];
              muxOutConnector[40] = fifoOut[38][3];
              muxOutConnector[41] = fifoOut[39][3];
              muxOutConnector[42] = fifoOut[40][3];
              muxOutConnector[43] = fifoOut[41][3];
              muxOutConnector[44] = fifoOut[42][3];
              muxOutConnector[45] = fifoOut[43][3];
              muxOutConnector[46] = fifoOut[44][3];
              muxOutConnector[47] = fifoOut[45][3];
              muxOutConnector[48] = fifoOut[46][3];
              muxOutConnector[49] = fifoOut[47][3];
              muxOutConnector[50] = fifoOut[48][3];
              muxOutConnector[51] = fifoOut[49][3];
         end
         14: begin
              muxOutConnector[0] = fifoOut[39][16];
              muxOutConnector[1] = fifoOut[40][16];
              muxOutConnector[2] = fifoOut[41][16];
              muxOutConnector[3] = fifoOut[42][16];
              muxOutConnector[4] = fifoOut[43][16];
              muxOutConnector[5] = fifoOut[44][16];
              muxOutConnector[6] = fifoOut[45][16];
              muxOutConnector[7] = fifoOut[46][16];
              muxOutConnector[8] = fifoOut[47][16];
              muxOutConnector[9] = fifoOut[48][16];
              muxOutConnector[10] = fifoOut[49][16];
              muxOutConnector[11] = fifoOut[50][16];
              muxOutConnector[12] = fifoOut[51][16];
              muxOutConnector[13] = fifoOut[26][15];
              muxOutConnector[14] = fifoOut[27][15];
              muxOutConnector[15] = fifoOut[28][15];
              muxOutConnector[16] = fifoOut[29][15];
              muxOutConnector[17] = fifoOut[30][15];
              muxOutConnector[18] = fifoOut[31][15];
              muxOutConnector[19] = fifoOut[32][15];
              muxOutConnector[20] = fifoOut[33][15];
              muxOutConnector[21] = fifoOut[34][15];
              muxOutConnector[22] = fifoOut[35][15];
              muxOutConnector[23] = fifoOut[36][15];
              muxOutConnector[24] = fifoOut[37][15];
              muxOutConnector[25] = fifoOut[38][15];
              muxOutConnector[26] = fifoOut[50][4];
              muxOutConnector[27] = fifoOut[51][4];
              muxOutConnector[28] = fifoOut[26][3];
              muxOutConnector[29] = fifoOut[27][3];
              muxOutConnector[30] = fifoOut[28][3];
              muxOutConnector[31] = fifoOut[29][3];
              muxOutConnector[32] = fifoOut[30][3];
              muxOutConnector[33] = fifoOut[31][3];
              muxOutConnector[34] = fifoOut[32][3];
              muxOutConnector[35] = fifoOut[33][3];
              muxOutConnector[36] = fifoOut[34][3];
              muxOutConnector[37] = fifoOut[35][3];
              muxOutConnector[38] = fifoOut[36][3];
              muxOutConnector[39] = fifoOut[37][3];
              muxOutConnector[40] = fifoOut[38][3];
              muxOutConnector[41] = fifoOut[39][3];
              muxOutConnector[42] = fifoOut[40][3];
              muxOutConnector[43] = fifoOut[41][3];
              muxOutConnector[44] = fifoOut[42][3];
              muxOutConnector[45] = fifoOut[43][3];
              muxOutConnector[46] = fifoOut[44][3];
              muxOutConnector[47] = fifoOut[45][3];
              muxOutConnector[48] = fifoOut[46][3];
              muxOutConnector[49] = fifoOut[47][3];
              muxOutConnector[50] = fifoOut[48][3];
              muxOutConnector[51] = fifoOut[49][3];
         end
         15: begin
              muxOutConnector[0] = fifoOut[39][16];
              muxOutConnector[1] = fifoOut[40][16];
              muxOutConnector[2] = fifoOut[41][16];
              muxOutConnector[3] = fifoOut[42][16];
              muxOutConnector[4] = fifoOut[43][16];
              muxOutConnector[5] = fifoOut[44][16];
              muxOutConnector[6] = fifoOut[45][16];
              muxOutConnector[7] = fifoOut[46][16];
              muxOutConnector[8] = fifoOut[47][16];
              muxOutConnector[9] = fifoOut[48][16];
              muxOutConnector[10] = fifoOut[49][16];
              muxOutConnector[11] = fifoOut[50][16];
              muxOutConnector[12] = fifoOut[51][16];
              muxOutConnector[13] = fifoOut[26][15];
              muxOutConnector[14] = fifoOut[27][15];
              muxOutConnector[15] = fifoOut[28][15];
              muxOutConnector[16] = fifoOut[29][15];
              muxOutConnector[17] = fifoOut[30][15];
              muxOutConnector[18] = fifoOut[31][15];
              muxOutConnector[19] = fifoOut[32][15];
              muxOutConnector[20] = fifoOut[33][15];
              muxOutConnector[21] = fifoOut[34][15];
              muxOutConnector[22] = fifoOut[35][15];
              muxOutConnector[23] = fifoOut[36][15];
              muxOutConnector[24] = fifoOut[37][15];
              muxOutConnector[25] = fifoOut[38][15];
              muxOutConnector[26] = fifoOut[50][4];
              muxOutConnector[27] = fifoOut[51][4];
              muxOutConnector[28] = fifoOut[26][3];
              muxOutConnector[29] = fifoOut[27][3];
              muxOutConnector[30] = fifoOut[28][3];
              muxOutConnector[31] = fifoOut[29][3];
              muxOutConnector[32] = fifoOut[30][3];
              muxOutConnector[33] = fifoOut[31][3];
              muxOutConnector[34] = fifoOut[32][3];
              muxOutConnector[35] = fifoOut[33][3];
              muxOutConnector[36] = fifoOut[34][3];
              muxOutConnector[37] = fifoOut[35][3];
              muxOutConnector[38] = fifoOut[36][3];
              muxOutConnector[39] = fifoOut[37][3];
              muxOutConnector[40] = fifoOut[38][3];
              muxOutConnector[41] = fifoOut[39][3];
              muxOutConnector[42] = fifoOut[40][3];
              muxOutConnector[43] = fifoOut[41][3];
              muxOutConnector[44] = fifoOut[42][3];
              muxOutConnector[45] = fifoOut[43][3];
              muxOutConnector[46] = fifoOut[44][3];
              muxOutConnector[47] = fifoOut[45][3];
              muxOutConnector[48] = fifoOut[46][3];
              muxOutConnector[49] = fifoOut[47][3];
              muxOutConnector[50] = fifoOut[48][3];
              muxOutConnector[51] = fifoOut[49][3];
         end
         16: begin
              muxOutConnector[0] = fifoOut[39][16];
              muxOutConnector[1] = fifoOut[40][16];
              muxOutConnector[2] = fifoOut[41][16];
              muxOutConnector[3] = fifoOut[42][16];
              muxOutConnector[4] = fifoOut[23][11];
              muxOutConnector[5] = fifoOut[24][11];
              muxOutConnector[6] = fifoOut[25][11];
              muxOutConnector[7] = fifoOut[0][10];
              muxOutConnector[8] = fifoOut[1][10];
              muxOutConnector[9] = fifoOut[2][10];
              muxOutConnector[10] = fifoOut[3][10];
              muxOutConnector[11] = fifoOut[4][10];
              muxOutConnector[12] = fifoOut[5][10];
              muxOutConnector[13] = fifoOut[6][10];
              muxOutConnector[14] = fifoOut[7][10];
              muxOutConnector[15] = fifoOut[8][10];
              muxOutConnector[16] = fifoOut[9][10];
              muxOutConnector[17] = fifoOut[10][10];
              muxOutConnector[18] = fifoOut[11][10];
              muxOutConnector[19] = fifoOut[12][10];
              muxOutConnector[20] = fifoOut[13][10];
              muxOutConnector[21] = fifoOut[14][10];
              muxOutConnector[22] = fifoOut[15][10];
              muxOutConnector[23] = fifoOut[16][10];
              muxOutConnector[24] = fifoOut[17][10];
              muxOutConnector[25] = fifoOut[18][10];
              muxOutConnector[26] = fifoOut[50][4];
              muxOutConnector[27] = fifoOut[51][4];
              muxOutConnector[28] = fifoOut[26][3];
              muxOutConnector[29] = fifoOut[27][3];
              muxOutConnector[30] = fifoOut[28][3];
              muxOutConnector[31] = fifoOut[29][3];
              muxOutConnector[32] = fifoOut[30][3];
              muxOutConnector[33] = fifoOut[31][3];
              muxOutConnector[34] = fifoOut[32][3];
              muxOutConnector[35] = fifoOut[33][3];
              muxOutConnector[36] = fifoOut[34][3];
              muxOutConnector[37] = fifoOut[35][3];
              muxOutConnector[38] = fifoOut[36][3];
              muxOutConnector[39] = fifoOut[37][3];
              muxOutConnector[40] = fifoOut[38][3];
              muxOutConnector[41] = fifoOut[39][3];
              muxOutConnector[42] = fifoOut[40][3];
              muxOutConnector[43] = fifoOut[41][3];
              muxOutConnector[44] = fifoOut[42][3];
              muxOutConnector[45] = fifoOut[43][3];
              muxOutConnector[46] = fifoOut[44][3];
              muxOutConnector[47] = fifoOut[45][3];
              muxOutConnector[48] = fifoOut[46][3];
              muxOutConnector[49] = fifoOut[47][3];
              muxOutConnector[50] = fifoOut[48][3];
              muxOutConnector[51] = fifoOut[49][3];
         end
         17: begin
              muxOutConnector[0] = fifoOut[19][11];
              muxOutConnector[1] = fifoOut[20][11];
              muxOutConnector[2] = fifoOut[21][11];
              muxOutConnector[3] = fifoOut[22][11];
              muxOutConnector[4] = fifoOut[23][11];
              muxOutConnector[5] = fifoOut[24][11];
              muxOutConnector[6] = fifoOut[25][11];
              muxOutConnector[7] = fifoOut[0][10];
              muxOutConnector[8] = fifoOut[1][10];
              muxOutConnector[9] = fifoOut[2][10];
              muxOutConnector[10] = fifoOut[3][10];
              muxOutConnector[11] = fifoOut[4][10];
              muxOutConnector[12] = fifoOut[5][10];
              muxOutConnector[13] = fifoOut[6][10];
              muxOutConnector[14] = fifoOut[7][10];
              muxOutConnector[15] = fifoOut[8][10];
              muxOutConnector[16] = fifoOut[9][10];
              muxOutConnector[17] = fifoOut[10][10];
              muxOutConnector[18] = fifoOut[11][10];
              muxOutConnector[19] = fifoOut[12][10];
              muxOutConnector[20] = fifoOut[13][10];
              muxOutConnector[21] = fifoOut[14][10];
              muxOutConnector[22] = fifoOut[15][10];
              muxOutConnector[23] = fifoOut[16][10];
              muxOutConnector[24] = fifoOut[17][10];
              muxOutConnector[25] = fifoOut[18][10];
              muxOutConnector[26] = fifoOut[50][4];
              muxOutConnector[27] = fifoOut[51][4];
              muxOutConnector[28] = fifoOut[26][3];
              muxOutConnector[29] = fifoOut[27][3];
              muxOutConnector[30] = fifoOut[28][3];
              muxOutConnector[31] = fifoOut[29][3];
              muxOutConnector[32] = fifoOut[30][3];
              muxOutConnector[33] = fifoOut[31][3];
              muxOutConnector[34] = fifoOut[32][3];
              muxOutConnector[35] = fifoOut[33][3];
              muxOutConnector[36] = fifoOut[34][3];
              muxOutConnector[37] = fifoOut[35][3];
              muxOutConnector[38] = fifoOut[36][3];
              muxOutConnector[39] = fifoOut[37][3];
              muxOutConnector[40] = fifoOut[38][3];
              muxOutConnector[41] = fifoOut[39][3];
              muxOutConnector[42] = fifoOut[40][3];
              muxOutConnector[43] = fifoOut[41][3];
              muxOutConnector[44] = fifoOut[42][3];
              muxOutConnector[45] = fifoOut[43][3];
              muxOutConnector[46] = fifoOut[44][3];
              muxOutConnector[47] = fifoOut[45][3];
              muxOutConnector[48] = fifoOut[46][3];
              muxOutConnector[49] = fifoOut[47][3];
              muxOutConnector[50] = fifoOut[48][3];
              muxOutConnector[51] = fifoOut[49][3];
         end
         18: begin
              muxOutConnector[0] = fifoOut[19][11];
              muxOutConnector[1] = fifoOut[20][11];
              muxOutConnector[2] = fifoOut[21][11];
              muxOutConnector[3] = fifoOut[22][11];
              muxOutConnector[4] = fifoOut[23][11];
              muxOutConnector[5] = fifoOut[24][11];
              muxOutConnector[6] = fifoOut[25][11];
              muxOutConnector[7] = fifoOut[0][10];
              muxOutConnector[8] = fifoOut[1][10];
              muxOutConnector[9] = fifoOut[2][10];
              muxOutConnector[10] = fifoOut[3][10];
              muxOutConnector[11] = fifoOut[4][10];
              muxOutConnector[12] = fifoOut[5][10];
              muxOutConnector[13] = fifoOut[6][10];
              muxOutConnector[14] = fifoOut[7][10];
              muxOutConnector[15] = fifoOut[8][10];
              muxOutConnector[16] = fifoOut[9][10];
              muxOutConnector[17] = fifoOut[10][10];
              muxOutConnector[18] = fifoOut[11][10];
              muxOutConnector[19] = fifoOut[12][10];
              muxOutConnector[20] = fifoOut[13][10];
              muxOutConnector[21] = fifoOut[14][10];
              muxOutConnector[22] = fifoOut[15][10];
              muxOutConnector[23] = fifoOut[16][10];
              muxOutConnector[24] = fifoOut[17][10];
              muxOutConnector[25] = fifoOut[18][10];
              muxOutConnector[26] = fifoOut[50][4];
              muxOutConnector[27] = fifoOut[51][4];
              muxOutConnector[28] = fifoOut[26][3];
              muxOutConnector[29] = fifoOut[27][3];
              muxOutConnector[30] = fifoOut[28][3];
              muxOutConnector[31] = fifoOut[29][3];
              muxOutConnector[32] = fifoOut[30][3];
              muxOutConnector[33] = fifoOut[31][3];
              muxOutConnector[34] = fifoOut[32][3];
              muxOutConnector[35] = fifoOut[33][3];
              muxOutConnector[36] = fifoOut[34][3];
              muxOutConnector[37] = fifoOut[35][3];
              muxOutConnector[38] = fifoOut[36][3];
              muxOutConnector[39] = fifoOut[37][3];
              muxOutConnector[40] = fifoOut[38][3];
              muxOutConnector[41] = fifoOut[39][3];
              muxOutConnector[42] = fifoOut[40][3];
              muxOutConnector[43] = fifoOut[41][3];
              muxOutConnector[44] = fifoOut[42][3];
              muxOutConnector[45] = fifoOut[43][3];
              muxOutConnector[46] = fifoOut[44][3];
              muxOutConnector[47] = fifoOut[45][3];
              muxOutConnector[48] = fifoOut[46][3];
              muxOutConnector[49] = fifoOut[47][3];
              muxOutConnector[50] = fifoOut[48][3];
              muxOutConnector[51] = fifoOut[49][3];
         end
         19: begin
              muxOutConnector[0] = fifoOut[19][11];
              muxOutConnector[1] = fifoOut[20][11];
              muxOutConnector[2] = fifoOut[21][11];
              muxOutConnector[3] = fifoOut[22][11];
              muxOutConnector[4] = fifoOut[23][11];
              muxOutConnector[5] = fifoOut[24][11];
              muxOutConnector[6] = fifoOut[25][11];
              muxOutConnector[7] = fifoOut[0][10];
              muxOutConnector[8] = fifoOut[1][10];
              muxOutConnector[9] = fifoOut[2][10];
              muxOutConnector[10] = fifoOut[3][10];
              muxOutConnector[11] = fifoOut[4][10];
              muxOutConnector[12] = fifoOut[5][10];
              muxOutConnector[13] = fifoOut[6][10];
              muxOutConnector[14] = fifoOut[7][10];
              muxOutConnector[15] = fifoOut[8][10];
              muxOutConnector[16] = fifoOut[9][10];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[50][4];
              muxOutConnector[27] = fifoOut[51][4];
              muxOutConnector[28] = fifoOut[26][3];
              muxOutConnector[29] = fifoOut[27][3];
              muxOutConnector[30] = fifoOut[28][3];
              muxOutConnector[31] = fifoOut[29][3];
              muxOutConnector[32] = fifoOut[30][3];
              muxOutConnector[33] = fifoOut[31][3];
              muxOutConnector[34] = fifoOut[32][3];
              muxOutConnector[35] = fifoOut[33][3];
              muxOutConnector[36] = fifoOut[34][3];
              muxOutConnector[37] = fifoOut[35][3];
              muxOutConnector[38] = fifoOut[36][3];
              muxOutConnector[39] = fifoOut[37][3];
              muxOutConnector[40] = fifoOut[38][3];
              muxOutConnector[41] = fifoOut[39][3];
              muxOutConnector[42] = fifoOut[40][3];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
         end
         default: begin
               for(i=0;i<muxOutSymbols;i=i+1)begin
                muxOutConnector[i] = 0;
              end
         end
//hgjhgbuiguigbigbgbgbui
         endcase
    end
endcase
             end
        endmodule