`timescale 1ns / 1ps
module LMem1To0_511_circ1_yesshift_nounload_scripted(
        muxOut,
        ly0In,
        wr_en,
        feedback_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 14;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

input feedback_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        if(feedback_en) begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= fifoOut[i][c-1];
         end
        end
        else begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= ly0InConnector[i];
         end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[3][4];
              muxOutConnector[1] = fifoOut[4][4];
              muxOutConnector[2] = fifoOut[5][4];
              muxOutConnector[3] = fifoOut[6][4];
              muxOutConnector[4] = fifoOut[7][4];
              muxOutConnector[5] = fifoOut[8][4];
              muxOutConnector[6] = fifoOut[9][4];
              muxOutConnector[7] = fifoOut[10][4];
              muxOutConnector[8] = fifoOut[11][4];
              muxOutConnector[9] = fifoOut[12][4];
              muxOutConnector[10] = fifoOut[13][4];
              muxOutConnector[11] = fifoOut[14][4];
              muxOutConnector[12] = fifoOut[15][4];
              muxOutConnector[13] = fifoOut[16][4];
              muxOutConnector[14] = fifoOut[17][4];
              muxOutConnector[15] = fifoOut[18][4];
              muxOutConnector[16] = fifoOut[19][4];
              muxOutConnector[17] = fifoOut[20][4];
              muxOutConnector[18] = fifoOut[21][4];
              muxOutConnector[19] = fifoOut[22][4];
              muxOutConnector[20] = fifoOut[23][4];
              muxOutConnector[21] = fifoOut[24][4];
              muxOutConnector[22] = fifoOut[25][4];
              muxOutConnector[23] = fifoOut[0][3];
              muxOutConnector[24] = fifoOut[1][3];
              muxOutConnector[25] = fifoOut[2][3];
              muxOutConnector[26] = fifoOut[43][9];
              muxOutConnector[27] = fifoOut[44][9];
              muxOutConnector[28] = fifoOut[45][9];
              muxOutConnector[29] = fifoOut[46][9];
              muxOutConnector[30] = fifoOut[47][9];
              muxOutConnector[31] = fifoOut[48][9];
              muxOutConnector[32] = fifoOut[49][9];
              muxOutConnector[33] = fifoOut[50][9];
              muxOutConnector[34] = fifoOut[51][9];
              muxOutConnector[35] = fifoOut[26][8];
              muxOutConnector[36] = fifoOut[27][8];
              muxOutConnector[37] = fifoOut[28][8];
              muxOutConnector[38] = fifoOut[29][8];
              muxOutConnector[39] = fifoOut[30][8];
              muxOutConnector[40] = fifoOut[31][8];
              muxOutConnector[41] = fifoOut[32][8];
              muxOutConnector[42] = fifoOut[33][8];
              muxOutConnector[43] = fifoOut[34][8];
              muxOutConnector[44] = fifoOut[35][8];
              muxOutConnector[45] = fifoOut[36][8];
              muxOutConnector[46] = fifoOut[37][8];
              muxOutConnector[47] = fifoOut[38][8];
              muxOutConnector[48] = fifoOut[39][8];
              muxOutConnector[49] = fifoOut[40][8];
              muxOutConnector[50] = fifoOut[41][8];
              muxOutConnector[51] = fifoOut[42][8];
       end
       1: begin
              muxOutConnector[0] = fifoOut[3][4];
              muxOutConnector[1] = fifoOut[4][4];
              muxOutConnector[2] = fifoOut[5][4];
              muxOutConnector[3] = fifoOut[6][4];
              muxOutConnector[4] = fifoOut[7][4];
              muxOutConnector[5] = fifoOut[8][4];
              muxOutConnector[6] = fifoOut[9][4];
              muxOutConnector[7] = fifoOut[10][4];
              muxOutConnector[8] = fifoOut[11][4];
              muxOutConnector[9] = fifoOut[12][4];
              muxOutConnector[10] = fifoOut[13][4];
              muxOutConnector[11] = fifoOut[14][4];
              muxOutConnector[12] = fifoOut[15][4];
              muxOutConnector[13] = fifoOut[16][4];
              muxOutConnector[14] = fifoOut[17][4];
              muxOutConnector[15] = fifoOut[18][4];
              muxOutConnector[16] = fifoOut[19][4];
              muxOutConnector[17] = fifoOut[20][4];
              muxOutConnector[18] = fifoOut[21][4];
              muxOutConnector[19] = fifoOut[22][4];
              muxOutConnector[20] = fifoOut[23][4];
              muxOutConnector[21] = fifoOut[24][4];
              muxOutConnector[22] = fifoOut[25][4];
              muxOutConnector[23] = fifoOut[0][3];
              muxOutConnector[24] = fifoOut[1][3];
              muxOutConnector[25] = fifoOut[2][3];
              muxOutConnector[26] = fifoOut[43][9];
              muxOutConnector[27] = fifoOut[44][9];
              muxOutConnector[28] = fifoOut[45][9];
              muxOutConnector[29] = fifoOut[46][9];
              muxOutConnector[30] = fifoOut[47][9];
              muxOutConnector[31] = fifoOut[48][9];
              muxOutConnector[32] = fifoOut[49][9];
              muxOutConnector[33] = fifoOut[50][9];
              muxOutConnector[34] = fifoOut[51][9];
              muxOutConnector[35] = fifoOut[26][8];
              muxOutConnector[36] = fifoOut[27][8];
              muxOutConnector[37] = fifoOut[28][8];
              muxOutConnector[38] = fifoOut[29][8];
              muxOutConnector[39] = fifoOut[30][8];
              muxOutConnector[40] = fifoOut[31][8];
              muxOutConnector[41] = fifoOut[32][8];
              muxOutConnector[42] = fifoOut[33][8];
              muxOutConnector[43] = fifoOut[34][8];
              muxOutConnector[44] = fifoOut[35][8];
              muxOutConnector[45] = fifoOut[36][8];
              muxOutConnector[46] = fifoOut[37][8];
              muxOutConnector[47] = fifoOut[38][8];
              muxOutConnector[48] = fifoOut[39][8];
              muxOutConnector[49] = fifoOut[40][8];
              muxOutConnector[50] = fifoOut[41][8];
              muxOutConnector[51] = fifoOut[42][8];
       end
       2: begin
              muxOutConnector[0] = fifoOut[3][4];
              muxOutConnector[1] = fifoOut[4][4];
              muxOutConnector[2] = fifoOut[5][4];
              muxOutConnector[3] = fifoOut[6][4];
              muxOutConnector[4] = fifoOut[7][4];
              muxOutConnector[5] = fifoOut[8][4];
              muxOutConnector[6] = fifoOut[9][4];
              muxOutConnector[7] = fifoOut[10][4];
              muxOutConnector[8] = fifoOut[11][4];
              muxOutConnector[9] = fifoOut[12][4];
              muxOutConnector[10] = fifoOut[13][4];
              muxOutConnector[11] = fifoOut[14][4];
              muxOutConnector[12] = fifoOut[15][4];
              muxOutConnector[13] = fifoOut[16][4];
              muxOutConnector[14] = fifoOut[17][4];
              muxOutConnector[15] = fifoOut[18][4];
              muxOutConnector[16] = fifoOut[19][4];
              muxOutConnector[17] = fifoOut[20][4];
              muxOutConnector[18] = fifoOut[21][4];
              muxOutConnector[19] = fifoOut[22][4];
              muxOutConnector[20] = fifoOut[23][4];
              muxOutConnector[21] = fifoOut[24][4];
              muxOutConnector[22] = fifoOut[25][4];
              muxOutConnector[23] = fifoOut[0][3];
              muxOutConnector[24] = fifoOut[1][3];
              muxOutConnector[25] = fifoOut[2][3];
              muxOutConnector[26] = fifoOut[43][9];
              muxOutConnector[27] = fifoOut[44][9];
              muxOutConnector[28] = fifoOut[45][9];
              muxOutConnector[29] = fifoOut[46][9];
              muxOutConnector[30] = fifoOut[47][9];
              muxOutConnector[31] = fifoOut[48][9];
              muxOutConnector[32] = fifoOut[49][9];
              muxOutConnector[33] = fifoOut[50][9];
              muxOutConnector[34] = fifoOut[51][9];
              muxOutConnector[35] = fifoOut[26][8];
              muxOutConnector[36] = fifoOut[27][8];
              muxOutConnector[37] = fifoOut[28][8];
              muxOutConnector[38] = fifoOut[29][8];
              muxOutConnector[39] = fifoOut[30][8];
              muxOutConnector[40] = fifoOut[31][8];
              muxOutConnector[41] = fifoOut[32][8];
              muxOutConnector[42] = fifoOut[33][8];
              muxOutConnector[43] = fifoOut[34][8];
              muxOutConnector[44] = fifoOut[35][8];
              muxOutConnector[45] = fifoOut[36][8];
              muxOutConnector[46] = fifoOut[37][8];
              muxOutConnector[47] = fifoOut[38][8];
              muxOutConnector[48] = fifoOut[39][8];
              muxOutConnector[49] = fifoOut[40][8];
              muxOutConnector[50] = fifoOut[41][8];
              muxOutConnector[51] = fifoOut[42][8];
       end
       3: begin
              muxOutConnector[0] = fifoOut[3][4];
              muxOutConnector[1] = fifoOut[4][4];
              muxOutConnector[2] = fifoOut[5][4];
              muxOutConnector[3] = fifoOut[6][4];
              muxOutConnector[4] = fifoOut[7][4];
              muxOutConnector[5] = fifoOut[8][4];
              muxOutConnector[6] = fifoOut[9][4];
              muxOutConnector[7] = fifoOut[10][4];
              muxOutConnector[8] = fifoOut[11][4];
              muxOutConnector[9] = fifoOut[12][4];
              muxOutConnector[10] = fifoOut[13][4];
              muxOutConnector[11] = fifoOut[14][4];
              muxOutConnector[12] = fifoOut[15][4];
              muxOutConnector[13] = fifoOut[16][4];
              muxOutConnector[14] = fifoOut[17][4];
              muxOutConnector[15] = fifoOut[18][4];
              muxOutConnector[16] = fifoOut[19][4];
              muxOutConnector[17] = fifoOut[20][4];
              muxOutConnector[18] = fifoOut[21][4];
              muxOutConnector[19] = fifoOut[22][4];
              muxOutConnector[20] = fifoOut[23][4];
              muxOutConnector[21] = fifoOut[24][4];
              muxOutConnector[22] = fifoOut[25][4];
              muxOutConnector[23] = fifoOut[0][3];
              muxOutConnector[24] = fifoOut[1][3];
              muxOutConnector[25] = fifoOut[2][3];
              muxOutConnector[26] = fifoOut[43][9];
              muxOutConnector[27] = fifoOut[44][9];
              muxOutConnector[28] = fifoOut[45][9];
              muxOutConnector[29] = fifoOut[46][9];
              muxOutConnector[30] = fifoOut[47][9];
              muxOutConnector[31] = fifoOut[48][9];
              muxOutConnector[32] = fifoOut[49][9];
              muxOutConnector[33] = fifoOut[50][9];
              muxOutConnector[34] = fifoOut[51][9];
              muxOutConnector[35] = fifoOut[26][8];
              muxOutConnector[36] = fifoOut[27][8];
              muxOutConnector[37] = fifoOut[28][8];
              muxOutConnector[38] = fifoOut[29][8];
              muxOutConnector[39] = fifoOut[30][8];
              muxOutConnector[40] = fifoOut[31][8];
              muxOutConnector[41] = fifoOut[32][8];
              muxOutConnector[42] = fifoOut[33][8];
              muxOutConnector[43] = fifoOut[34][8];
              muxOutConnector[44] = fifoOut[35][8];
              muxOutConnector[45] = fifoOut[36][8];
              muxOutConnector[46] = fifoOut[37][8];
              muxOutConnector[47] = fifoOut[38][8];
              muxOutConnector[48] = fifoOut[39][8];
              muxOutConnector[49] = fifoOut[40][8];
              muxOutConnector[50] = fifoOut[41][8];
              muxOutConnector[51] = fifoOut[42][8];
       end
       4: begin
              muxOutConnector[0] = fifoOut[3][4];
              muxOutConnector[1] = fifoOut[4][4];
              muxOutConnector[2] = fifoOut[5][4];
              muxOutConnector[3] = fifoOut[6][4];
              muxOutConnector[4] = fifoOut[7][4];
              muxOutConnector[5] = fifoOut[8][4];
              muxOutConnector[6] = fifoOut[9][4];
              muxOutConnector[7] = fifoOut[10][4];
              muxOutConnector[8] = fifoOut[11][4];
              muxOutConnector[9] = fifoOut[12][4];
              muxOutConnector[10] = fifoOut[13][4];
              muxOutConnector[11] = fifoOut[14][4];
              muxOutConnector[12] = fifoOut[15][4];
              muxOutConnector[13] = fifoOut[16][4];
              muxOutConnector[14] = fifoOut[38][3];
              muxOutConnector[15] = fifoOut[39][3];
              muxOutConnector[16] = fifoOut[40][3];
              muxOutConnector[17] = fifoOut[41][3];
              muxOutConnector[18] = fifoOut[42][3];
              muxOutConnector[19] = fifoOut[43][3];
              muxOutConnector[20] = fifoOut[44][3];
              muxOutConnector[21] = fifoOut[45][3];
              muxOutConnector[22] = fifoOut[46][3];
              muxOutConnector[23] = fifoOut[47][3];
              muxOutConnector[24] = fifoOut[48][3];
              muxOutConnector[25] = fifoOut[49][3];
              muxOutConnector[26] = fifoOut[43][9];
              muxOutConnector[27] = fifoOut[44][9];
              muxOutConnector[28] = fifoOut[45][9];
              muxOutConnector[29] = fifoOut[46][9];
              muxOutConnector[30] = fifoOut[47][9];
              muxOutConnector[31] = fifoOut[48][9];
              muxOutConnector[32] = fifoOut[49][9];
              muxOutConnector[33] = fifoOut[50][9];
              muxOutConnector[34] = fifoOut[51][9];
              muxOutConnector[35] = fifoOut[26][8];
              muxOutConnector[36] = fifoOut[27][8];
              muxOutConnector[37] = fifoOut[28][8];
              muxOutConnector[38] = fifoOut[29][8];
              muxOutConnector[39] = fifoOut[30][8];
              muxOutConnector[40] = fifoOut[31][8];
              muxOutConnector[41] = fifoOut[32][8];
              muxOutConnector[42] = fifoOut[33][8];
              muxOutConnector[43] = fifoOut[34][8];
              muxOutConnector[44] = fifoOut[35][8];
              muxOutConnector[45] = fifoOut[36][8];
              muxOutConnector[46] = fifoOut[37][8];
              muxOutConnector[47] = fifoOut[38][8];
              muxOutConnector[48] = fifoOut[39][8];
              muxOutConnector[49] = fifoOut[40][8];
              muxOutConnector[50] = fifoOut[41][8];
              muxOutConnector[51] = fifoOut[42][8];
       end
       5: begin
              muxOutConnector[0] = fifoOut[50][4];
              muxOutConnector[1] = fifoOut[51][4];
              muxOutConnector[2] = fifoOut[26][3];
              muxOutConnector[3] = fifoOut[27][3];
              muxOutConnector[4] = fifoOut[28][3];
              muxOutConnector[5] = fifoOut[29][3];
              muxOutConnector[6] = fifoOut[30][3];
              muxOutConnector[7] = fifoOut[31][3];
              muxOutConnector[8] = fifoOut[32][3];
              muxOutConnector[9] = fifoOut[33][3];
              muxOutConnector[10] = fifoOut[34][3];
              muxOutConnector[11] = fifoOut[35][3];
              muxOutConnector[12] = fifoOut[36][3];
              muxOutConnector[13] = fifoOut[37][3];
              muxOutConnector[14] = fifoOut[38][3];
              muxOutConnector[15] = fifoOut[39][3];
              muxOutConnector[16] = fifoOut[40][3];
              muxOutConnector[17] = fifoOut[41][3];
              muxOutConnector[18] = fifoOut[42][3];
              muxOutConnector[19] = fifoOut[43][3];
              muxOutConnector[20] = fifoOut[44][3];
              muxOutConnector[21] = fifoOut[45][3];
              muxOutConnector[22] = fifoOut[46][3];
              muxOutConnector[23] = fifoOut[47][3];
              muxOutConnector[24] = fifoOut[48][3];
              muxOutConnector[25] = fifoOut[49][3];
              muxOutConnector[26] = fifoOut[43][9];
              muxOutConnector[27] = fifoOut[44][9];
              muxOutConnector[28] = fifoOut[45][9];
              muxOutConnector[29] = fifoOut[46][9];
              muxOutConnector[30] = fifoOut[47][9];
              muxOutConnector[31] = fifoOut[48][9];
              muxOutConnector[32] = fifoOut[49][9];
              muxOutConnector[33] = fifoOut[50][9];
              muxOutConnector[34] = fifoOut[51][9];
              muxOutConnector[35] = fifoOut[26][8];
              muxOutConnector[36] = fifoOut[27][8];
              muxOutConnector[37] = fifoOut[28][8];
              muxOutConnector[38] = fifoOut[29][8];
              muxOutConnector[39] = fifoOut[30][8];
              muxOutConnector[40] = fifoOut[31][8];
              muxOutConnector[41] = fifoOut[32][8];
              muxOutConnector[42] = fifoOut[33][8];
              muxOutConnector[43] = fifoOut[34][8];
              muxOutConnector[44] = fifoOut[35][8];
              muxOutConnector[45] = fifoOut[36][8];
              muxOutConnector[46] = fifoOut[37][8];
              muxOutConnector[47] = fifoOut[38][8];
              muxOutConnector[48] = fifoOut[39][8];
              muxOutConnector[49] = fifoOut[40][8];
              muxOutConnector[50] = fifoOut[41][8];
              muxOutConnector[51] = fifoOut[42][8];
       end
       6: begin
              muxOutConnector[0] = fifoOut[50][4];
              muxOutConnector[1] = fifoOut[51][4];
              muxOutConnector[2] = fifoOut[26][3];
              muxOutConnector[3] = fifoOut[27][3];
              muxOutConnector[4] = fifoOut[28][3];
              muxOutConnector[5] = fifoOut[29][3];
              muxOutConnector[6] = fifoOut[30][3];
              muxOutConnector[7] = fifoOut[31][3];
              muxOutConnector[8] = fifoOut[32][3];
              muxOutConnector[9] = fifoOut[33][3];
              muxOutConnector[10] = fifoOut[34][3];
              muxOutConnector[11] = fifoOut[35][3];
              muxOutConnector[12] = fifoOut[36][3];
              muxOutConnector[13] = fifoOut[37][3];
              muxOutConnector[14] = fifoOut[38][3];
              muxOutConnector[15] = fifoOut[39][3];
              muxOutConnector[16] = fifoOut[40][3];
              muxOutConnector[17] = fifoOut[41][3];
              muxOutConnector[18] = fifoOut[42][3];
              muxOutConnector[19] = fifoOut[43][3];
              muxOutConnector[20] = fifoOut[44][3];
              muxOutConnector[21] = fifoOut[45][3];
              muxOutConnector[22] = fifoOut[46][3];
              muxOutConnector[23] = fifoOut[47][3];
              muxOutConnector[24] = fifoOut[48][3];
              muxOutConnector[25] = fifoOut[49][3];
              muxOutConnector[26] = fifoOut[43][9];
              muxOutConnector[27] = fifoOut[44][9];
              muxOutConnector[28] = fifoOut[45][9];
              muxOutConnector[29] = fifoOut[46][9];
              muxOutConnector[30] = fifoOut[47][9];
              muxOutConnector[31] = fifoOut[48][9];
              muxOutConnector[32] = fifoOut[49][9];
              muxOutConnector[33] = fifoOut[50][9];
              muxOutConnector[34] = fifoOut[51][9];
              muxOutConnector[35] = fifoOut[26][8];
              muxOutConnector[36] = fifoOut[27][8];
              muxOutConnector[37] = fifoOut[28][8];
              muxOutConnector[38] = fifoOut[29][8];
              muxOutConnector[39] = fifoOut[30][8];
              muxOutConnector[40] = fifoOut[31][8];
              muxOutConnector[41] = fifoOut[32][8];
              muxOutConnector[42] = fifoOut[33][8];
              muxOutConnector[43] = fifoOut[34][8];
              muxOutConnector[44] = fifoOut[35][8];
              muxOutConnector[45] = fifoOut[36][8];
              muxOutConnector[46] = fifoOut[37][8];
              muxOutConnector[47] = fifoOut[38][8];
              muxOutConnector[48] = fifoOut[39][8];
              muxOutConnector[49] = fifoOut[40][8];
              muxOutConnector[50] = fifoOut[41][8];
              muxOutConnector[51] = fifoOut[42][8];
       end
       7: begin
              muxOutConnector[0] = fifoOut[50][4];
              muxOutConnector[1] = fifoOut[51][4];
              muxOutConnector[2] = fifoOut[26][3];
              muxOutConnector[3] = fifoOut[27][3];
              muxOutConnector[4] = fifoOut[28][3];
              muxOutConnector[5] = fifoOut[29][3];
              muxOutConnector[6] = fifoOut[30][3];
              muxOutConnector[7] = fifoOut[31][3];
              muxOutConnector[8] = fifoOut[32][3];
              muxOutConnector[9] = fifoOut[33][3];
              muxOutConnector[10] = fifoOut[34][3];
              muxOutConnector[11] = fifoOut[35][3];
              muxOutConnector[12] = fifoOut[36][3];
              muxOutConnector[13] = fifoOut[37][3];
              muxOutConnector[14] = fifoOut[38][3];
              muxOutConnector[15] = fifoOut[39][3];
              muxOutConnector[16] = fifoOut[40][3];
              muxOutConnector[17] = fifoOut[41][3];
              muxOutConnector[18] = fifoOut[42][3];
              muxOutConnector[19] = fifoOut[43][3];
              muxOutConnector[20] = fifoOut[44][3];
              muxOutConnector[21] = fifoOut[45][3];
              muxOutConnector[22] = fifoOut[46][3];
              muxOutConnector[23] = fifoOut[47][3];
              muxOutConnector[24] = fifoOut[48][3];
              muxOutConnector[25] = fifoOut[49][3];
              muxOutConnector[26] = fifoOut[43][9];
              muxOutConnector[27] = fifoOut[44][9];
              muxOutConnector[28] = fifoOut[45][9];
              muxOutConnector[29] = fifoOut[46][9];
              muxOutConnector[30] = fifoOut[47][9];
              muxOutConnector[31] = fifoOut[48][9];
              muxOutConnector[32] = fifoOut[49][9];
              muxOutConnector[33] = fifoOut[50][9];
              muxOutConnector[34] = fifoOut[51][9];
              muxOutConnector[35] = fifoOut[26][8];
              muxOutConnector[36] = fifoOut[27][8];
              muxOutConnector[37] = fifoOut[28][8];
              muxOutConnector[38] = fifoOut[29][8];
              muxOutConnector[39] = fifoOut[30][8];
              muxOutConnector[40] = fifoOut[31][8];
              muxOutConnector[41] = fifoOut[32][8];
              muxOutConnector[42] = fifoOut[33][8];
              muxOutConnector[43] = fifoOut[34][8];
              muxOutConnector[44] = fifoOut[35][8];
              muxOutConnector[45] = fifoOut[36][8];
              muxOutConnector[46] = fifoOut[37][8];
              muxOutConnector[47] = fifoOut[38][8];
              muxOutConnector[48] = fifoOut[39][8];
              muxOutConnector[49] = fifoOut[40][8];
              muxOutConnector[50] = fifoOut[41][8];
              muxOutConnector[51] = fifoOut[42][8];
       end
       8: begin
              muxOutConnector[0] = fifoOut[50][4];
              muxOutConnector[1] = fifoOut[51][4];
              muxOutConnector[2] = fifoOut[26][3];
              muxOutConnector[3] = fifoOut[27][3];
              muxOutConnector[4] = fifoOut[28][3];
              muxOutConnector[5] = fifoOut[29][3];
              muxOutConnector[6] = fifoOut[30][3];
              muxOutConnector[7] = fifoOut[31][3];
              muxOutConnector[8] = fifoOut[32][3];
              muxOutConnector[9] = fifoOut[33][3];
              muxOutConnector[10] = fifoOut[34][3];
              muxOutConnector[11] = fifoOut[35][3];
              muxOutConnector[12] = fifoOut[36][3];
              muxOutConnector[13] = fifoOut[37][3];
              muxOutConnector[14] = fifoOut[38][3];
              muxOutConnector[15] = fifoOut[39][3];
              muxOutConnector[16] = fifoOut[40][3];
              muxOutConnector[17] = fifoOut[41][3];
              muxOutConnector[18] = fifoOut[42][3];
              muxOutConnector[19] = fifoOut[43][3];
              muxOutConnector[20] = fifoOut[44][3];
              muxOutConnector[21] = fifoOut[45][3];
              muxOutConnector[22] = fifoOut[46][3];
              muxOutConnector[23] = fifoOut[47][3];
              muxOutConnector[24] = fifoOut[48][3];
              muxOutConnector[25] = fifoOut[49][3];
              muxOutConnector[26] = fifoOut[43][9];
              muxOutConnector[27] = fifoOut[44][9];
              muxOutConnector[28] = fifoOut[45][9];
              muxOutConnector[29] = fifoOut[46][9];
              muxOutConnector[30] = fifoOut[47][9];
              muxOutConnector[31] = fifoOut[48][9];
              muxOutConnector[32] = fifoOut[49][9];
              muxOutConnector[33] = fifoOut[50][9];
              muxOutConnector[34] = fifoOut[51][9];
              muxOutConnector[35] = fifoOut[26][8];
              muxOutConnector[36] = fifoOut[27][8];
              muxOutConnector[37] = fifoOut[28][8];
              muxOutConnector[38] = fifoOut[29][8];
              muxOutConnector[39] = fifoOut[30][8];
              muxOutConnector[40] = fifoOut[31][8];
              muxOutConnector[41] = fifoOut[32][8];
              muxOutConnector[42] = fifoOut[33][8];
              muxOutConnector[43] = fifoOut[34][8];
              muxOutConnector[44] = fifoOut[35][8];
              muxOutConnector[45] = fifoOut[36][8];
              muxOutConnector[46] = fifoOut[37][8];
              muxOutConnector[47] = fifoOut[38][8];
              muxOutConnector[48] = fifoOut[39][8];
              muxOutConnector[49] = fifoOut[40][8];
              muxOutConnector[50] = fifoOut[41][8];
              muxOutConnector[51] = fifoOut[42][8];
       end
       9: begin
              muxOutConnector[0] = fifoOut[50][4];
              muxOutConnector[1] = fifoOut[51][4];
              muxOutConnector[2] = fifoOut[26][3];
              muxOutConnector[3] = fifoOut[27][3];
              muxOutConnector[4] = fifoOut[28][3];
              muxOutConnector[5] = fifoOut[29][3];
              muxOutConnector[6] = fifoOut[30][3];
              muxOutConnector[7] = fifoOut[31][3];
              muxOutConnector[8] = fifoOut[32][3];
              muxOutConnector[9] = fifoOut[33][3];
              muxOutConnector[10] = fifoOut[34][3];
              muxOutConnector[11] = fifoOut[35][3];
              muxOutConnector[12] = fifoOut[36][3];
              muxOutConnector[13] = fifoOut[37][3];
              muxOutConnector[14] = fifoOut[38][3];
              muxOutConnector[15] = fifoOut[39][3];
              muxOutConnector[16] = fifoOut[40][3];
              muxOutConnector[17] = fifoOut[41][3];
              muxOutConnector[18] = fifoOut[42][3];
              muxOutConnector[19] = fifoOut[43][3];
              muxOutConnector[20] = fifoOut[44][3];
              muxOutConnector[21] = fifoOut[45][3];
              muxOutConnector[22] = fifoOut[46][3];
              muxOutConnector[23] = fifoOut[47][3];
              muxOutConnector[24] = fifoOut[48][3];
              muxOutConnector[25] = fifoOut[49][3];
              muxOutConnector[26] = fifoOut[5][1];
              muxOutConnector[27] = fifoOut[6][1];
              muxOutConnector[28] = fifoOut[7][1];
              muxOutConnector[29] = fifoOut[8][1];
              muxOutConnector[30] = fifoOut[9][1];
              muxOutConnector[31] = fifoOut[10][1];
              muxOutConnector[32] = fifoOut[11][1];
              muxOutConnector[33] = fifoOut[12][1];
              muxOutConnector[34] = fifoOut[13][1];
              muxOutConnector[35] = fifoOut[14][1];
              muxOutConnector[36] = fifoOut[15][1];
              muxOutConnector[37] = fifoOut[16][1];
              muxOutConnector[38] = fifoOut[17][1];
              muxOutConnector[39] = fifoOut[18][1];
              muxOutConnector[40] = fifoOut[19][1];
              muxOutConnector[41] = fifoOut[20][1];
              muxOutConnector[42] = fifoOut[21][1];
              muxOutConnector[43] = fifoOut[22][1];
              muxOutConnector[44] = fifoOut[23][1];
              muxOutConnector[45] = fifoOut[24][1];
              muxOutConnector[46] = fifoOut[25][1];
              muxOutConnector[47] = fifoOut[0][0];
              muxOutConnector[48] = fifoOut[1][0];
              muxOutConnector[49] = fifoOut[2][0];
              muxOutConnector[50] = fifoOut[3][0];
              muxOutConnector[51] = fifoOut[4][0];
       end
       10: begin
              muxOutConnector[0] = fifoOut[50][4];
              muxOutConnector[1] = fifoOut[51][4];
              muxOutConnector[2] = fifoOut[26][3];
              muxOutConnector[3] = fifoOut[27][3];
              muxOutConnector[4] = fifoOut[28][3];
              muxOutConnector[5] = fifoOut[29][3];
              muxOutConnector[6] = fifoOut[30][3];
              muxOutConnector[7] = fifoOut[31][3];
              muxOutConnector[8] = fifoOut[32][3];
              muxOutConnector[9] = fifoOut[33][3];
              muxOutConnector[10] = fifoOut[34][3];
              muxOutConnector[11] = fifoOut[35][3];
              muxOutConnector[12] = fifoOut[36][3];
              muxOutConnector[13] = fifoOut[37][3];
              muxOutConnector[14] = fifoOut[0][9];
              muxOutConnector[15] = fifoOut[1][9];
              muxOutConnector[16] = fifoOut[2][9];
              muxOutConnector[17] = fifoOut[3][9];
              muxOutConnector[18] = fifoOut[4][9];
              muxOutConnector[19] = fifoOut[5][9];
              muxOutConnector[20] = fifoOut[6][9];
              muxOutConnector[21] = fifoOut[7][9];
              muxOutConnector[22] = fifoOut[8][9];
              muxOutConnector[23] = fifoOut[9][9];
              muxOutConnector[24] = fifoOut[10][9];
              muxOutConnector[25] = fifoOut[11][9];
              muxOutConnector[26] = fifoOut[5][1];
              muxOutConnector[27] = fifoOut[6][1];
              muxOutConnector[28] = fifoOut[7][1];
              muxOutConnector[29] = fifoOut[8][1];
              muxOutConnector[30] = fifoOut[9][1];
              muxOutConnector[31] = fifoOut[10][1];
              muxOutConnector[32] = fifoOut[11][1];
              muxOutConnector[33] = fifoOut[12][1];
              muxOutConnector[34] = fifoOut[13][1];
              muxOutConnector[35] = fifoOut[14][1];
              muxOutConnector[36] = fifoOut[15][1];
              muxOutConnector[37] = fifoOut[16][1];
              muxOutConnector[38] = fifoOut[17][1];
              muxOutConnector[39] = fifoOut[18][1];
              muxOutConnector[40] = fifoOut[19][1];
              muxOutConnector[41] = fifoOut[20][1];
              muxOutConnector[42] = fifoOut[21][1];
              muxOutConnector[43] = fifoOut[22][1];
              muxOutConnector[44] = fifoOut[23][1];
              muxOutConnector[45] = fifoOut[24][1];
              muxOutConnector[46] = fifoOut[25][1];
              muxOutConnector[47] = fifoOut[0][0];
              muxOutConnector[48] = fifoOut[1][0];
              muxOutConnector[49] = fifoOut[2][0];
              muxOutConnector[50] = fifoOut[3][0];
              muxOutConnector[51] = fifoOut[4][0];
       end
       11: begin
              muxOutConnector[0] = fifoOut[12][10];
              muxOutConnector[1] = fifoOut[13][10];
              muxOutConnector[2] = fifoOut[14][10];
              muxOutConnector[3] = fifoOut[15][10];
              muxOutConnector[4] = fifoOut[16][10];
              muxOutConnector[5] = fifoOut[17][10];
              muxOutConnector[6] = fifoOut[18][10];
              muxOutConnector[7] = fifoOut[19][10];
              muxOutConnector[8] = fifoOut[20][10];
              muxOutConnector[9] = fifoOut[21][10];
              muxOutConnector[10] = fifoOut[22][10];
              muxOutConnector[11] = fifoOut[23][10];
              muxOutConnector[12] = fifoOut[24][10];
              muxOutConnector[13] = fifoOut[25][10];
              muxOutConnector[14] = fifoOut[0][9];
              muxOutConnector[15] = fifoOut[1][9];
              muxOutConnector[16] = fifoOut[2][9];
              muxOutConnector[17] = fifoOut[3][9];
              muxOutConnector[18] = fifoOut[4][9];
              muxOutConnector[19] = fifoOut[5][9];
              muxOutConnector[20] = fifoOut[6][9];
              muxOutConnector[21] = fifoOut[7][9];
              muxOutConnector[22] = fifoOut[8][9];
              muxOutConnector[23] = fifoOut[9][9];
              muxOutConnector[24] = fifoOut[10][9];
              muxOutConnector[25] = fifoOut[11][9];
              muxOutConnector[26] = fifoOut[5][1];
              muxOutConnector[27] = fifoOut[6][1];
              muxOutConnector[28] = fifoOut[7][1];
              muxOutConnector[29] = fifoOut[8][1];
              muxOutConnector[30] = fifoOut[9][1];
              muxOutConnector[31] = fifoOut[10][1];
              muxOutConnector[32] = fifoOut[11][1];
              muxOutConnector[33] = fifoOut[12][1];
              muxOutConnector[34] = fifoOut[13][1];
              muxOutConnector[35] = fifoOut[14][1];
              muxOutConnector[36] = fifoOut[15][1];
              muxOutConnector[37] = fifoOut[16][1];
              muxOutConnector[38] = fifoOut[17][1];
              muxOutConnector[39] = fifoOut[18][1];
              muxOutConnector[40] = fifoOut[19][1];
              muxOutConnector[41] = fifoOut[20][1];
              muxOutConnector[42] = fifoOut[21][1];
              muxOutConnector[43] = fifoOut[22][1];
              muxOutConnector[44] = fifoOut[23][1];
              muxOutConnector[45] = fifoOut[24][1];
              muxOutConnector[46] = fifoOut[25][1];
              muxOutConnector[47] = fifoOut[0][0];
              muxOutConnector[48] = fifoOut[1][0];
              muxOutConnector[49] = fifoOut[2][0];
              muxOutConnector[50] = fifoOut[3][0];
              muxOutConnector[51] = fifoOut[4][0];
       end
       12: begin
              muxOutConnector[0] = fifoOut[12][10];
              muxOutConnector[1] = fifoOut[13][10];
              muxOutConnector[2] = fifoOut[14][10];
              muxOutConnector[3] = fifoOut[15][10];
              muxOutConnector[4] = fifoOut[16][10];
              muxOutConnector[5] = fifoOut[17][10];
              muxOutConnector[6] = fifoOut[18][10];
              muxOutConnector[7] = fifoOut[19][10];
              muxOutConnector[8] = fifoOut[20][10];
              muxOutConnector[9] = fifoOut[21][10];
              muxOutConnector[10] = fifoOut[22][10];
              muxOutConnector[11] = fifoOut[23][10];
              muxOutConnector[12] = fifoOut[24][10];
              muxOutConnector[13] = fifoOut[25][10];
              muxOutConnector[14] = fifoOut[0][9];
              muxOutConnector[15] = fifoOut[1][9];
              muxOutConnector[16] = fifoOut[2][9];
              muxOutConnector[17] = fifoOut[3][9];
              muxOutConnector[18] = fifoOut[4][9];
              muxOutConnector[19] = fifoOut[5][9];
              muxOutConnector[20] = fifoOut[6][9];
              muxOutConnector[21] = fifoOut[7][9];
              muxOutConnector[22] = fifoOut[8][9];
              muxOutConnector[23] = fifoOut[9][9];
              muxOutConnector[24] = fifoOut[10][9];
              muxOutConnector[25] = fifoOut[11][9];
              muxOutConnector[26] = fifoOut[5][1];
              muxOutConnector[27] = fifoOut[6][1];
              muxOutConnector[28] = fifoOut[7][1];
              muxOutConnector[29] = fifoOut[8][1];
              muxOutConnector[30] = fifoOut[9][1];
              muxOutConnector[31] = fifoOut[10][1];
              muxOutConnector[32] = fifoOut[11][1];
              muxOutConnector[33] = fifoOut[12][1];
              muxOutConnector[34] = fifoOut[13][1];
              muxOutConnector[35] = fifoOut[14][1];
              muxOutConnector[36] = fifoOut[15][1];
              muxOutConnector[37] = fifoOut[16][1];
              muxOutConnector[38] = fifoOut[17][1];
              muxOutConnector[39] = fifoOut[18][1];
              muxOutConnector[40] = fifoOut[19][1];
              muxOutConnector[41] = fifoOut[20][1];
              muxOutConnector[42] = fifoOut[21][1];
              muxOutConnector[43] = fifoOut[22][1];
              muxOutConnector[44] = fifoOut[23][1];
              muxOutConnector[45] = fifoOut[24][1];
              muxOutConnector[46] = fifoOut[25][1];
              muxOutConnector[47] = fifoOut[0][0];
              muxOutConnector[48] = fifoOut[1][0];
              muxOutConnector[49] = fifoOut[2][0];
              muxOutConnector[50] = fifoOut[3][0];
              muxOutConnector[51] = fifoOut[4][0];
       end
       13: begin
              muxOutConnector[0] = fifoOut[12][10];
              muxOutConnector[1] = fifoOut[13][10];
              muxOutConnector[2] = fifoOut[14][10];
              muxOutConnector[3] = fifoOut[15][10];
              muxOutConnector[4] = fifoOut[16][10];
              muxOutConnector[5] = fifoOut[17][10];
              muxOutConnector[6] = fifoOut[18][10];
              muxOutConnector[7] = fifoOut[19][10];
              muxOutConnector[8] = fifoOut[20][10];
              muxOutConnector[9] = fifoOut[21][10];
              muxOutConnector[10] = fifoOut[22][10];
              muxOutConnector[11] = fifoOut[23][10];
              muxOutConnector[12] = fifoOut[24][10];
              muxOutConnector[13] = fifoOut[25][10];
              muxOutConnector[14] = fifoOut[0][9];
              muxOutConnector[15] = fifoOut[1][9];
              muxOutConnector[16] = fifoOut[2][9];
              muxOutConnector[17] = fifoOut[3][9];
              muxOutConnector[18] = fifoOut[4][9];
              muxOutConnector[19] = fifoOut[5][9];
              muxOutConnector[20] = fifoOut[6][9];
              muxOutConnector[21] = fifoOut[7][9];
              muxOutConnector[22] = fifoOut[8][9];
              muxOutConnector[23] = fifoOut[9][9];
              muxOutConnector[24] = fifoOut[10][9];
              muxOutConnector[25] = fifoOut[11][9];
              muxOutConnector[26] = fifoOut[5][1];
              muxOutConnector[27] = fifoOut[6][1];
              muxOutConnector[28] = fifoOut[7][1];
              muxOutConnector[29] = fifoOut[8][1];
              muxOutConnector[30] = fifoOut[9][1];
              muxOutConnector[31] = fifoOut[10][1];
              muxOutConnector[32] = fifoOut[11][1];
              muxOutConnector[33] = fifoOut[12][1];
              muxOutConnector[34] = fifoOut[13][1];
              muxOutConnector[35] = fifoOut[14][1];
              muxOutConnector[36] = fifoOut[15][1];
              muxOutConnector[37] = fifoOut[16][1];
              muxOutConnector[38] = fifoOut[17][1];
              muxOutConnector[39] = fifoOut[18][1];
              muxOutConnector[40] = fifoOut[19][1];
              muxOutConnector[41] = fifoOut[20][1];
              muxOutConnector[42] = fifoOut[21][1];
              muxOutConnector[43] = fifoOut[22][1];
              muxOutConnector[44] = fifoOut[23][1];
              muxOutConnector[45] = fifoOut[24][1];
              muxOutConnector[46] = fifoOut[25][1];
              muxOutConnector[47] = fifoOut[0][0];
              muxOutConnector[48] = fifoOut[1][0];
              muxOutConnector[49] = fifoOut[2][0];
              muxOutConnector[50] = fifoOut[3][0];
              muxOutConnector[51] = fifoOut[4][0];
       end
       14: begin
              muxOutConnector[0] = fifoOut[12][10];
              muxOutConnector[1] = fifoOut[13][10];
              muxOutConnector[2] = fifoOut[14][10];
              muxOutConnector[3] = fifoOut[15][10];
              muxOutConnector[4] = fifoOut[16][10];
              muxOutConnector[5] = fifoOut[17][10];
              muxOutConnector[6] = fifoOut[18][10];
              muxOutConnector[7] = fifoOut[19][10];
              muxOutConnector[8] = fifoOut[20][10];
              muxOutConnector[9] = fifoOut[21][10];
              muxOutConnector[10] = fifoOut[22][10];
              muxOutConnector[11] = fifoOut[23][10];
              muxOutConnector[12] = fifoOut[24][10];
              muxOutConnector[13] = fifoOut[25][10];
              muxOutConnector[14] = fifoOut[0][9];
              muxOutConnector[15] = fifoOut[1][9];
              muxOutConnector[16] = fifoOut[2][9];
              muxOutConnector[17] = fifoOut[3][9];
              muxOutConnector[18] = fifoOut[4][9];
              muxOutConnector[19] = fifoOut[5][9];
              muxOutConnector[20] = fifoOut[6][9];
              muxOutConnector[21] = fifoOut[7][9];
              muxOutConnector[22] = fifoOut[8][9];
              muxOutConnector[23] = fifoOut[9][9];
              muxOutConnector[24] = fifoOut[10][9];
              muxOutConnector[25] = fifoOut[11][9];
              muxOutConnector[26] = fifoOut[5][1];
              muxOutConnector[27] = fifoOut[6][1];
              muxOutConnector[28] = fifoOut[7][1];
              muxOutConnector[29] = fifoOut[8][1];
              muxOutConnector[30] = fifoOut[9][1];
              muxOutConnector[31] = fifoOut[10][1];
              muxOutConnector[32] = fifoOut[11][1];
              muxOutConnector[33] = fifoOut[12][1];
              muxOutConnector[34] = fifoOut[13][1];
              muxOutConnector[35] = fifoOut[14][1];
              muxOutConnector[36] = fifoOut[15][1];
              muxOutConnector[37] = fifoOut[16][1];
              muxOutConnector[38] = fifoOut[17][1];
              muxOutConnector[39] = fifoOut[18][1];
              muxOutConnector[40] = fifoOut[19][1];
              muxOutConnector[41] = fifoOut[20][1];
              muxOutConnector[42] = fifoOut[21][1];
              muxOutConnector[43] = fifoOut[22][1];
              muxOutConnector[44] = fifoOut[23][1];
              muxOutConnector[45] = fifoOut[24][1];
              muxOutConnector[46] = fifoOut[25][1];
              muxOutConnector[47] = fifoOut[0][0];
              muxOutConnector[48] = fifoOut[1][0];
              muxOutConnector[49] = fifoOut[2][0];
              muxOutConnector[50] = fifoOut[3][0];
              muxOutConnector[51] = fifoOut[4][0];
       end
       15: begin
              muxOutConnector[0] = fifoOut[12][10];
              muxOutConnector[1] = fifoOut[13][10];
              muxOutConnector[2] = fifoOut[14][10];
              muxOutConnector[3] = fifoOut[15][10];
              muxOutConnector[4] = fifoOut[16][10];
              muxOutConnector[5] = fifoOut[17][10];
              muxOutConnector[6] = fifoOut[18][10];
              muxOutConnector[7] = fifoOut[19][10];
              muxOutConnector[8] = fifoOut[20][10];
              muxOutConnector[9] = fifoOut[21][10];
              muxOutConnector[10] = fifoOut[22][10];
              muxOutConnector[11] = fifoOut[23][10];
              muxOutConnector[12] = fifoOut[24][10];
              muxOutConnector[13] = fifoOut[25][10];
              muxOutConnector[14] = fifoOut[0][9];
              muxOutConnector[15] = fifoOut[1][9];
              muxOutConnector[16] = fifoOut[2][9];
              muxOutConnector[17] = fifoOut[3][9];
              muxOutConnector[18] = fifoOut[4][9];
              muxOutConnector[19] = fifoOut[5][9];
              muxOutConnector[20] = fifoOut[6][9];
              muxOutConnector[21] = fifoOut[7][9];
              muxOutConnector[22] = fifoOut[8][9];
              muxOutConnector[23] = fifoOut[9][9];
              muxOutConnector[24] = fifoOut[10][9];
              muxOutConnector[25] = fifoOut[11][9];
              muxOutConnector[26] = fifoOut[5][1];
              muxOutConnector[27] = fifoOut[6][1];
              muxOutConnector[28] = fifoOut[7][1];
              muxOutConnector[29] = fifoOut[8][1];
              muxOutConnector[30] = fifoOut[9][1];
              muxOutConnector[31] = fifoOut[10][1];
              muxOutConnector[32] = fifoOut[11][1];
              muxOutConnector[33] = fifoOut[12][1];
              muxOutConnector[34] = fifoOut[13][1];
              muxOutConnector[35] = fifoOut[14][1];
              muxOutConnector[36] = fifoOut[15][1];
              muxOutConnector[37] = fifoOut[16][1];
              muxOutConnector[38] = fifoOut[38][0];
              muxOutConnector[39] = fifoOut[39][0];
              muxOutConnector[40] = fifoOut[40][0];
              muxOutConnector[41] = fifoOut[41][0];
              muxOutConnector[42] = fifoOut[42][0];
              muxOutConnector[43] = fifoOut[43][0];
              muxOutConnector[44] = fifoOut[44][0];
              muxOutConnector[45] = fifoOut[45][0];
              muxOutConnector[46] = fifoOut[46][0];
              muxOutConnector[47] = fifoOut[47][0];
              muxOutConnector[48] = fifoOut[48][0];
              muxOutConnector[49] = fifoOut[49][0];
              muxOutConnector[50] = fifoOut[50][0];
              muxOutConnector[51] = fifoOut[51][0];
       end
       16: begin
              muxOutConnector[0] = fifoOut[12][10];
              muxOutConnector[1] = fifoOut[13][10];
              muxOutConnector[2] = fifoOut[14][10];
              muxOutConnector[3] = fifoOut[15][10];
              muxOutConnector[4] = fifoOut[16][10];
              muxOutConnector[5] = fifoOut[17][10];
              muxOutConnector[6] = fifoOut[18][10];
              muxOutConnector[7] = fifoOut[19][10];
              muxOutConnector[8] = fifoOut[20][10];
              muxOutConnector[9] = fifoOut[21][10];
              muxOutConnector[10] = fifoOut[22][10];
              muxOutConnector[11] = fifoOut[23][10];
              muxOutConnector[12] = fifoOut[24][10];
              muxOutConnector[13] = fifoOut[25][10];
              muxOutConnector[14] = fifoOut[0][9];
              muxOutConnector[15] = fifoOut[1][9];
              muxOutConnector[16] = fifoOut[2][9];
              muxOutConnector[17] = fifoOut[3][9];
              muxOutConnector[18] = fifoOut[4][9];
              muxOutConnector[19] = fifoOut[5][9];
              muxOutConnector[20] = fifoOut[6][9];
              muxOutConnector[21] = fifoOut[7][9];
              muxOutConnector[22] = fifoOut[8][9];
              muxOutConnector[23] = fifoOut[9][9];
              muxOutConnector[24] = fifoOut[10][9];
              muxOutConnector[25] = fifoOut[11][9];
              muxOutConnector[26] = fifoOut[26][0];
              muxOutConnector[27] = fifoOut[27][0];
              muxOutConnector[28] = fifoOut[28][0];
              muxOutConnector[29] = fifoOut[29][0];
              muxOutConnector[30] = fifoOut[30][0];
              muxOutConnector[31] = fifoOut[31][0];
              muxOutConnector[32] = fifoOut[32][0];
              muxOutConnector[33] = fifoOut[33][0];
              muxOutConnector[34] = fifoOut[34][0];
              muxOutConnector[35] = fifoOut[35][0];
              muxOutConnector[36] = fifoOut[36][0];
              muxOutConnector[37] = fifoOut[37][0];
              muxOutConnector[38] = fifoOut[38][0];
              muxOutConnector[39] = fifoOut[39][0];
              muxOutConnector[40] = fifoOut[40][0];
              muxOutConnector[41] = fifoOut[41][0];
              muxOutConnector[42] = fifoOut[42][0];
              muxOutConnector[43] = fifoOut[43][0];
              muxOutConnector[44] = fifoOut[44][0];
              muxOutConnector[45] = fifoOut[45][0];
              muxOutConnector[46] = fifoOut[46][0];
              muxOutConnector[47] = fifoOut[47][0];
              muxOutConnector[48] = fifoOut[48][0];
              muxOutConnector[49] = fifoOut[49][0];
              muxOutConnector[50] = fifoOut[50][0];
              muxOutConnector[51] = fifoOut[51][0];
       end
       17: begin
              muxOutConnector[0] = fifoOut[12][10];
              muxOutConnector[1] = fifoOut[13][10];
              muxOutConnector[2] = fifoOut[14][10];
              muxOutConnector[3] = fifoOut[15][10];
              muxOutConnector[4] = fifoOut[16][10];
              muxOutConnector[5] = fifoOut[17][10];
              muxOutConnector[6] = fifoOut[18][10];
              muxOutConnector[7] = fifoOut[19][10];
              muxOutConnector[8] = fifoOut[20][10];
              muxOutConnector[9] = fifoOut[21][10];
              muxOutConnector[10] = fifoOut[22][10];
              muxOutConnector[11] = fifoOut[23][10];
              muxOutConnector[12] = fifoOut[24][10];
              muxOutConnector[13] = fifoOut[25][10];
              muxOutConnector[14] = fifoOut[0][9];
              muxOutConnector[15] = fifoOut[1][9];
              muxOutConnector[16] = fifoOut[2][9];
              muxOutConnector[17] = fifoOut[3][9];
              muxOutConnector[18] = fifoOut[4][9];
              muxOutConnector[19] = fifoOut[5][9];
              muxOutConnector[20] = fifoOut[6][9];
              muxOutConnector[21] = fifoOut[7][9];
              muxOutConnector[22] = fifoOut[8][9];
              muxOutConnector[23] = fifoOut[9][9];
              muxOutConnector[24] = fifoOut[10][9];
              muxOutConnector[25] = fifoOut[11][9];
              muxOutConnector[26] = fifoOut[26][0];
              muxOutConnector[27] = fifoOut[27][0];
              muxOutConnector[28] = fifoOut[28][0];
              muxOutConnector[29] = fifoOut[29][0];
              muxOutConnector[30] = fifoOut[30][0];
              muxOutConnector[31] = fifoOut[31][0];
              muxOutConnector[32] = fifoOut[32][0];
              muxOutConnector[33] = fifoOut[33][0];
              muxOutConnector[34] = fifoOut[34][0];
              muxOutConnector[35] = fifoOut[35][0];
              muxOutConnector[36] = fifoOut[36][0];
              muxOutConnector[37] = fifoOut[37][0];
              muxOutConnector[38] = fifoOut[38][0];
              muxOutConnector[39] = fifoOut[39][0];
              muxOutConnector[40] = fifoOut[40][0];
              muxOutConnector[41] = fifoOut[41][0];
              muxOutConnector[42] = fifoOut[42][0];
              muxOutConnector[43] = fifoOut[43][0];
              muxOutConnector[44] = fifoOut[44][0];
              muxOutConnector[45] = fifoOut[45][0];
              muxOutConnector[46] = fifoOut[46][0];
              muxOutConnector[47] = fifoOut[47][0];
              muxOutConnector[48] = fifoOut[48][0];
              muxOutConnector[49] = fifoOut[49][0];
              muxOutConnector[50] = fifoOut[50][0];
              muxOutConnector[51] = fifoOut[51][0];
       end
       18: begin
              muxOutConnector[0] = fifoOut[12][10];
              muxOutConnector[1] = fifoOut[13][10];
              muxOutConnector[2] = fifoOut[14][10];
              muxOutConnector[3] = fifoOut[15][10];
              muxOutConnector[4] = fifoOut[16][10];
              muxOutConnector[5] = fifoOut[17][10];
              muxOutConnector[6] = fifoOut[18][10];
              muxOutConnector[7] = fifoOut[19][10];
              muxOutConnector[8] = fifoOut[20][10];
              muxOutConnector[9] = fifoOut[21][10];
              muxOutConnector[10] = fifoOut[22][10];
              muxOutConnector[11] = fifoOut[23][10];
              muxOutConnector[12] = fifoOut[24][10];
              muxOutConnector[13] = fifoOut[25][10];
              muxOutConnector[14] = fifoOut[0][9];
              muxOutConnector[15] = fifoOut[1][9];
              muxOutConnector[16] = fifoOut[2][9];
              muxOutConnector[17] = fifoOut[3][9];
              muxOutConnector[18] = fifoOut[4][9];
              muxOutConnector[19] = fifoOut[5][9];
              muxOutConnector[20] = fifoOut[6][9];
              muxOutConnector[21] = fifoOut[7][9];
              muxOutConnector[22] = fifoOut[8][9];
              muxOutConnector[23] = fifoOut[9][9];
              muxOutConnector[24] = fifoOut[10][9];
              muxOutConnector[25] = fifoOut[11][9];
              muxOutConnector[26] = fifoOut[26][0];
              muxOutConnector[27] = fifoOut[27][0];
              muxOutConnector[28] = fifoOut[28][0];
              muxOutConnector[29] = fifoOut[29][0];
              muxOutConnector[30] = fifoOut[30][0];
              muxOutConnector[31] = fifoOut[31][0];
              muxOutConnector[32] = fifoOut[32][0];
              muxOutConnector[33] = fifoOut[33][0];
              muxOutConnector[34] = fifoOut[34][0];
              muxOutConnector[35] = fifoOut[35][0];
              muxOutConnector[36] = fifoOut[36][0];
              muxOutConnector[37] = fifoOut[37][0];
              muxOutConnector[38] = fifoOut[38][0];
              muxOutConnector[39] = fifoOut[39][0];
              muxOutConnector[40] = fifoOut[40][0];
              muxOutConnector[41] = fifoOut[41][0];
              muxOutConnector[42] = fifoOut[42][0];
              muxOutConnector[43] = fifoOut[43][0];
              muxOutConnector[44] = fifoOut[44][0];
              muxOutConnector[45] = fifoOut[45][0];
              muxOutConnector[46] = fifoOut[46][0];
              muxOutConnector[47] = fifoOut[47][0];
              muxOutConnector[48] = fifoOut[48][0];
              muxOutConnector[49] = fifoOut[49][0];
              muxOutConnector[50] = fifoOut[50][0];
              muxOutConnector[51] = fifoOut[51][0];
       end
       19: begin
              muxOutConnector[0] = fifoOut[12][10];
              muxOutConnector[1] = fifoOut[13][10];
              muxOutConnector[2] = fifoOut[14][10];
              muxOutConnector[3] = fifoOut[15][10];
              muxOutConnector[4] = fifoOut[16][10];
              muxOutConnector[5] = fifoOut[17][10];
              muxOutConnector[6] = fifoOut[18][10];
              muxOutConnector[7] = fifoOut[19][10];
              muxOutConnector[8] = fifoOut[20][10];
              muxOutConnector[9] = fifoOut[21][10];
              muxOutConnector[10] = fifoOut[22][10];
              muxOutConnector[11] = fifoOut[23][10];
              muxOutConnector[12] = fifoOut[24][10];
              muxOutConnector[13] = fifoOut[25][10];
              muxOutConnector[14] = fifoOut[0][9];
              muxOutConnector[15] = fifoOut[1][9];
              muxOutConnector[16] = fifoOut[2][9];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[26][0];
              muxOutConnector[27] = fifoOut[27][0];
              muxOutConnector[28] = fifoOut[28][0];
              muxOutConnector[29] = fifoOut[29][0];
              muxOutConnector[30] = fifoOut[30][0];
              muxOutConnector[31] = fifoOut[31][0];
              muxOutConnector[32] = fifoOut[32][0];
              muxOutConnector[33] = fifoOut[33][0];
              muxOutConnector[34] = fifoOut[34][0];
              muxOutConnector[35] = fifoOut[35][0];
              muxOutConnector[36] = fifoOut[36][0];
              muxOutConnector[37] = fifoOut[37][0];
              muxOutConnector[38] = fifoOut[38][0];
              muxOutConnector[39] = fifoOut[39][0];
              muxOutConnector[40] = fifoOut[40][0];
              muxOutConnector[41] = fifoOut[41][0];
              muxOutConnector[42] = fifoOut[42][0];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
