`timescale 1ns / 1ps
module LMem1To0_511_circ5_yesshift_nounload_scripted(
        muxOut,
        ly0In,
        wr_en,
        feedback_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 13;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

input feedback_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        if(feedback_en) begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= fifoOut[i][c-1];
         end
        end
        else begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= ly0InConnector[i];
         end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[16][5];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[49][3];
              muxOutConnector[27] = fifoOut[50][3];
              muxOutConnector[28] = fifoOut[51][3];
              muxOutConnector[29] = fifoOut[26][2];
              muxOutConnector[30] = fifoOut[27][2];
              muxOutConnector[31] = fifoOut[28][2];
              muxOutConnector[32] = fifoOut[29][2];
              muxOutConnector[33] = fifoOut[30][2];
              muxOutConnector[34] = fifoOut[31][2];
              muxOutConnector[35] = fifoOut[32][2];
              muxOutConnector[36] = fifoOut[33][2];
              muxOutConnector[37] = fifoOut[34][2];
              muxOutConnector[38] = fifoOut[35][2];
              muxOutConnector[39] = fifoOut[36][2];
              muxOutConnector[40] = fifoOut[37][2];
              muxOutConnector[41] = fifoOut[38][2];
              muxOutConnector[42] = fifoOut[39][2];
              muxOutConnector[43] = fifoOut[40][2];
              muxOutConnector[44] = fifoOut[41][2];
              muxOutConnector[45] = fifoOut[42][2];
              muxOutConnector[46] = fifoOut[43][2];
              muxOutConnector[47] = fifoOut[44][2];
              muxOutConnector[48] = fifoOut[45][2];
              muxOutConnector[49] = fifoOut[46][2];
              muxOutConnector[50] = fifoOut[47][2];
              muxOutConnector[51] = fifoOut[48][2];
       end
       1: begin
              muxOutConnector[0] = fifoOut[16][5];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[49][3];
              muxOutConnector[27] = fifoOut[50][3];
              muxOutConnector[28] = fifoOut[51][3];
              muxOutConnector[29] = fifoOut[26][2];
              muxOutConnector[30] = fifoOut[27][2];
              muxOutConnector[31] = fifoOut[28][2];
              muxOutConnector[32] = fifoOut[29][2];
              muxOutConnector[33] = fifoOut[30][2];
              muxOutConnector[34] = fifoOut[31][2];
              muxOutConnector[35] = fifoOut[32][2];
              muxOutConnector[36] = fifoOut[33][2];
              muxOutConnector[37] = fifoOut[34][2];
              muxOutConnector[38] = fifoOut[35][2];
              muxOutConnector[39] = fifoOut[36][2];
              muxOutConnector[40] = fifoOut[37][2];
              muxOutConnector[41] = fifoOut[38][2];
              muxOutConnector[42] = fifoOut[39][2];
              muxOutConnector[43] = fifoOut[40][2];
              muxOutConnector[44] = fifoOut[41][2];
              muxOutConnector[45] = fifoOut[42][2];
              muxOutConnector[46] = fifoOut[43][2];
              muxOutConnector[47] = fifoOut[44][2];
              muxOutConnector[48] = fifoOut[45][2];
              muxOutConnector[49] = fifoOut[46][2];
              muxOutConnector[50] = fifoOut[47][2];
              muxOutConnector[51] = fifoOut[48][2];
       end
       2: begin
              muxOutConnector[0] = fifoOut[16][5];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[49][3];
              muxOutConnector[27] = fifoOut[50][3];
              muxOutConnector[28] = fifoOut[51][3];
              muxOutConnector[29] = fifoOut[26][2];
              muxOutConnector[30] = fifoOut[27][2];
              muxOutConnector[31] = fifoOut[28][2];
              muxOutConnector[32] = fifoOut[29][2];
              muxOutConnector[33] = fifoOut[30][2];
              muxOutConnector[34] = fifoOut[31][2];
              muxOutConnector[35] = fifoOut[32][2];
              muxOutConnector[36] = fifoOut[33][2];
              muxOutConnector[37] = fifoOut[34][2];
              muxOutConnector[38] = fifoOut[35][2];
              muxOutConnector[39] = fifoOut[36][2];
              muxOutConnector[40] = fifoOut[37][2];
              muxOutConnector[41] = fifoOut[38][2];
              muxOutConnector[42] = fifoOut[39][2];
              muxOutConnector[43] = fifoOut[40][2];
              muxOutConnector[44] = fifoOut[41][2];
              muxOutConnector[45] = fifoOut[42][2];
              muxOutConnector[46] = fifoOut[17][1];
              muxOutConnector[47] = fifoOut[18][1];
              muxOutConnector[48] = fifoOut[19][1];
              muxOutConnector[49] = fifoOut[20][1];
              muxOutConnector[50] = fifoOut[21][1];
              muxOutConnector[51] = fifoOut[22][1];
       end
       3: begin
              muxOutConnector[0] = fifoOut[16][5];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[23][2];
              muxOutConnector[27] = fifoOut[24][2];
              muxOutConnector[28] = fifoOut[25][2];
              muxOutConnector[29] = fifoOut[0][1];
              muxOutConnector[30] = fifoOut[1][1];
              muxOutConnector[31] = fifoOut[2][1];
              muxOutConnector[32] = fifoOut[3][1];
              muxOutConnector[33] = fifoOut[4][1];
              muxOutConnector[34] = fifoOut[5][1];
              muxOutConnector[35] = fifoOut[6][1];
              muxOutConnector[36] = fifoOut[7][1];
              muxOutConnector[37] = fifoOut[8][1];
              muxOutConnector[38] = fifoOut[9][1];
              muxOutConnector[39] = fifoOut[10][1];
              muxOutConnector[40] = fifoOut[11][1];
              muxOutConnector[41] = fifoOut[12][1];
              muxOutConnector[42] = fifoOut[13][1];
              muxOutConnector[43] = fifoOut[14][1];
              muxOutConnector[44] = fifoOut[15][1];
              muxOutConnector[45] = fifoOut[16][1];
              muxOutConnector[46] = fifoOut[17][1];
              muxOutConnector[47] = fifoOut[18][1];
              muxOutConnector[48] = fifoOut[19][1];
              muxOutConnector[49] = fifoOut[20][1];
              muxOutConnector[50] = fifoOut[21][1];
              muxOutConnector[51] = fifoOut[22][1];
       end
       4: begin
              muxOutConnector[0] = fifoOut[16][5];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[23][2];
              muxOutConnector[27] = fifoOut[24][2];
              muxOutConnector[28] = fifoOut[25][2];
              muxOutConnector[29] = fifoOut[0][1];
              muxOutConnector[30] = fifoOut[1][1];
              muxOutConnector[31] = fifoOut[2][1];
              muxOutConnector[32] = fifoOut[3][1];
              muxOutConnector[33] = fifoOut[4][1];
              muxOutConnector[34] = fifoOut[5][1];
              muxOutConnector[35] = fifoOut[6][1];
              muxOutConnector[36] = fifoOut[7][1];
              muxOutConnector[37] = fifoOut[8][1];
              muxOutConnector[38] = fifoOut[9][1];
              muxOutConnector[39] = fifoOut[10][1];
              muxOutConnector[40] = fifoOut[11][1];
              muxOutConnector[41] = fifoOut[12][1];
              muxOutConnector[42] = fifoOut[13][1];
              muxOutConnector[43] = fifoOut[14][1];
              muxOutConnector[44] = fifoOut[15][1];
              muxOutConnector[45] = fifoOut[16][1];
              muxOutConnector[46] = fifoOut[17][1];
              muxOutConnector[47] = fifoOut[18][1];
              muxOutConnector[48] = fifoOut[19][1];
              muxOutConnector[49] = fifoOut[20][1];
              muxOutConnector[50] = fifoOut[21][1];
              muxOutConnector[51] = fifoOut[22][1];
       end
       5: begin
              muxOutConnector[0] = fifoOut[16][5];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[23][2];
              muxOutConnector[27] = fifoOut[24][2];
              muxOutConnector[28] = fifoOut[25][2];
              muxOutConnector[29] = fifoOut[0][1];
              muxOutConnector[30] = fifoOut[1][1];
              muxOutConnector[31] = fifoOut[2][1];
              muxOutConnector[32] = fifoOut[3][1];
              muxOutConnector[33] = fifoOut[4][1];
              muxOutConnector[34] = fifoOut[5][1];
              muxOutConnector[35] = fifoOut[6][1];
              muxOutConnector[36] = fifoOut[7][1];
              muxOutConnector[37] = fifoOut[8][1];
              muxOutConnector[38] = fifoOut[9][1];
              muxOutConnector[39] = fifoOut[10][1];
              muxOutConnector[40] = fifoOut[11][1];
              muxOutConnector[41] = fifoOut[12][1];
              muxOutConnector[42] = fifoOut[13][1];
              muxOutConnector[43] = fifoOut[14][1];
              muxOutConnector[44] = fifoOut[15][1];
              muxOutConnector[45] = fifoOut[16][1];
              muxOutConnector[46] = fifoOut[17][1];
              muxOutConnector[47] = fifoOut[18][1];
              muxOutConnector[48] = fifoOut[19][1];
              muxOutConnector[49] = fifoOut[20][1];
              muxOutConnector[50] = fifoOut[21][1];
              muxOutConnector[51] = fifoOut[22][1];
       end
       6: begin
              muxOutConnector[0] = fifoOut[51][0];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[23][2];
              muxOutConnector[27] = fifoOut[24][2];
              muxOutConnector[28] = fifoOut[25][2];
              muxOutConnector[29] = fifoOut[0][1];
              muxOutConnector[30] = fifoOut[1][1];
              muxOutConnector[31] = fifoOut[2][1];
              muxOutConnector[32] = fifoOut[3][1];
              muxOutConnector[33] = fifoOut[4][1];
              muxOutConnector[34] = fifoOut[5][1];
              muxOutConnector[35] = fifoOut[6][1];
              muxOutConnector[36] = fifoOut[7][1];
              muxOutConnector[37] = fifoOut[8][1];
              muxOutConnector[38] = fifoOut[9][1];
              muxOutConnector[39] = fifoOut[10][1];
              muxOutConnector[40] = fifoOut[11][1];
              muxOutConnector[41] = fifoOut[12][1];
              muxOutConnector[42] = fifoOut[13][1];
              muxOutConnector[43] = fifoOut[14][1];
              muxOutConnector[44] = fifoOut[15][1];
              muxOutConnector[45] = fifoOut[16][1];
              muxOutConnector[46] = fifoOut[17][1];
              muxOutConnector[47] = fifoOut[18][1];
              muxOutConnector[48] = fifoOut[19][1];
              muxOutConnector[49] = fifoOut[20][1];
              muxOutConnector[50] = fifoOut[21][1];
              muxOutConnector[51] = fifoOut[22][1];
       end
       7: begin
              muxOutConnector[0] = fifoOut[51][0];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[23][2];
              muxOutConnector[27] = fifoOut[24][2];
              muxOutConnector[28] = fifoOut[25][2];
              muxOutConnector[29] = fifoOut[0][1];
              muxOutConnector[30] = fifoOut[1][1];
              muxOutConnector[31] = fifoOut[2][1];
              muxOutConnector[32] = fifoOut[3][1];
              muxOutConnector[33] = fifoOut[4][1];
              muxOutConnector[34] = fifoOut[5][1];
              muxOutConnector[35] = fifoOut[6][1];
              muxOutConnector[36] = fifoOut[7][1];
              muxOutConnector[37] = fifoOut[8][1];
              muxOutConnector[38] = fifoOut[9][1];
              muxOutConnector[39] = fifoOut[10][1];
              muxOutConnector[40] = fifoOut[11][1];
              muxOutConnector[41] = fifoOut[12][1];
              muxOutConnector[42] = fifoOut[13][1];
              muxOutConnector[43] = fifoOut[14][1];
              muxOutConnector[44] = fifoOut[15][1];
              muxOutConnector[45] = fifoOut[16][1];
              muxOutConnector[46] = fifoOut[17][1];
              muxOutConnector[47] = fifoOut[18][1];
              muxOutConnector[48] = fifoOut[19][1];
              muxOutConnector[49] = fifoOut[20][1];
              muxOutConnector[50] = fifoOut[21][1];
              muxOutConnector[51] = fifoOut[22][1];
       end
       8: begin
              muxOutConnector[0] = fifoOut[51][0];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[23][2];
              muxOutConnector[27] = fifoOut[24][2];
              muxOutConnector[28] = fifoOut[25][2];
              muxOutConnector[29] = fifoOut[0][1];
              muxOutConnector[30] = fifoOut[1][1];
              muxOutConnector[31] = fifoOut[2][1];
              muxOutConnector[32] = fifoOut[3][1];
              muxOutConnector[33] = fifoOut[4][1];
              muxOutConnector[34] = fifoOut[5][1];
              muxOutConnector[35] = fifoOut[6][1];
              muxOutConnector[36] = fifoOut[7][1];
              muxOutConnector[37] = fifoOut[8][1];
              muxOutConnector[38] = fifoOut[9][1];
              muxOutConnector[39] = fifoOut[10][1];
              muxOutConnector[40] = fifoOut[11][1];
              muxOutConnector[41] = fifoOut[12][1];
              muxOutConnector[42] = fifoOut[13][1];
              muxOutConnector[43] = fifoOut[14][1];
              muxOutConnector[44] = fifoOut[15][1];
              muxOutConnector[45] = fifoOut[16][1];
              muxOutConnector[46] = fifoOut[17][1];
              muxOutConnector[47] = fifoOut[18][1];
              muxOutConnector[48] = fifoOut[19][1];
              muxOutConnector[49] = fifoOut[20][1];
              muxOutConnector[50] = fifoOut[21][1];
              muxOutConnector[51] = fifoOut[22][1];
       end
       9: begin
              muxOutConnector[0] = fifoOut[51][0];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[23][2];
              muxOutConnector[27] = fifoOut[24][2];
              muxOutConnector[28] = fifoOut[25][2];
              muxOutConnector[29] = fifoOut[0][1];
              muxOutConnector[30] = fifoOut[1][1];
              muxOutConnector[31] = fifoOut[2][1];
              muxOutConnector[32] = fifoOut[3][1];
              muxOutConnector[33] = fifoOut[4][1];
              muxOutConnector[34] = fifoOut[5][1];
              muxOutConnector[35] = fifoOut[6][1];
              muxOutConnector[36] = fifoOut[7][1];
              muxOutConnector[37] = fifoOut[8][1];
              muxOutConnector[38] = fifoOut[9][1];
              muxOutConnector[39] = fifoOut[10][1];
              muxOutConnector[40] = fifoOut[11][1];
              muxOutConnector[41] = fifoOut[12][1];
              muxOutConnector[42] = fifoOut[13][1];
              muxOutConnector[43] = fifoOut[14][1];
              muxOutConnector[44] = fifoOut[15][1];
              muxOutConnector[45] = fifoOut[16][1];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       10: begin
              muxOutConnector[0] = fifoOut[51][0];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       11: begin
              muxOutConnector[0] = fifoOut[51][0];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[43][12];
              muxOutConnector[19] = fifoOut[44][12];
              muxOutConnector[20] = fifoOut[45][12];
              muxOutConnector[21] = fifoOut[46][12];
              muxOutConnector[22] = fifoOut[47][12];
              muxOutConnector[23] = fifoOut[48][12];
              muxOutConnector[24] = fifoOut[49][12];
              muxOutConnector[25] = fifoOut[50][12];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       12: begin
              muxOutConnector[0] = fifoOut[51][0];
              muxOutConnector[1] = fifoOut[26][12];
              muxOutConnector[2] = fifoOut[27][12];
              muxOutConnector[3] = fifoOut[28][12];
              muxOutConnector[4] = fifoOut[29][12];
              muxOutConnector[5] = fifoOut[30][12];
              muxOutConnector[6] = fifoOut[31][12];
              muxOutConnector[7] = fifoOut[32][12];
              muxOutConnector[8] = fifoOut[33][12];
              muxOutConnector[9] = fifoOut[34][12];
              muxOutConnector[10] = fifoOut[35][12];
              muxOutConnector[11] = fifoOut[36][12];
              muxOutConnector[12] = fifoOut[37][12];
              muxOutConnector[13] = fifoOut[38][12];
              muxOutConnector[14] = fifoOut[39][12];
              muxOutConnector[15] = fifoOut[40][12];
              muxOutConnector[16] = fifoOut[41][12];
              muxOutConnector[17] = fifoOut[42][12];
              muxOutConnector[18] = fifoOut[17][11];
              muxOutConnector[19] = fifoOut[18][11];
              muxOutConnector[20] = fifoOut[19][11];
              muxOutConnector[21] = fifoOut[20][11];
              muxOutConnector[22] = fifoOut[21][11];
              muxOutConnector[23] = fifoOut[22][11];
              muxOutConnector[24] = fifoOut[23][11];
              muxOutConnector[25] = fifoOut[24][11];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       13: begin
              muxOutConnector[0] = fifoOut[25][12];
              muxOutConnector[1] = fifoOut[0][11];
              muxOutConnector[2] = fifoOut[1][11];
              muxOutConnector[3] = fifoOut[2][11];
              muxOutConnector[4] = fifoOut[3][11];
              muxOutConnector[5] = fifoOut[4][11];
              muxOutConnector[6] = fifoOut[5][11];
              muxOutConnector[7] = fifoOut[6][11];
              muxOutConnector[8] = fifoOut[7][11];
              muxOutConnector[9] = fifoOut[8][11];
              muxOutConnector[10] = fifoOut[9][11];
              muxOutConnector[11] = fifoOut[10][11];
              muxOutConnector[12] = fifoOut[11][11];
              muxOutConnector[13] = fifoOut[12][11];
              muxOutConnector[14] = fifoOut[13][11];
              muxOutConnector[15] = fifoOut[14][11];
              muxOutConnector[16] = fifoOut[15][11];
              muxOutConnector[17] = fifoOut[16][11];
              muxOutConnector[18] = fifoOut[17][11];
              muxOutConnector[19] = fifoOut[18][11];
              muxOutConnector[20] = fifoOut[19][11];
              muxOutConnector[21] = fifoOut[20][11];
              muxOutConnector[22] = fifoOut[21][11];
              muxOutConnector[23] = fifoOut[22][11];
              muxOutConnector[24] = fifoOut[23][11];
              muxOutConnector[25] = fifoOut[24][11];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       14: begin
              muxOutConnector[0] = fifoOut[25][12];
              muxOutConnector[1] = fifoOut[0][11];
              muxOutConnector[2] = fifoOut[1][11];
              muxOutConnector[3] = fifoOut[2][11];
              muxOutConnector[4] = fifoOut[3][11];
              muxOutConnector[5] = fifoOut[4][11];
              muxOutConnector[6] = fifoOut[5][11];
              muxOutConnector[7] = fifoOut[6][11];
              muxOutConnector[8] = fifoOut[7][11];
              muxOutConnector[9] = fifoOut[8][11];
              muxOutConnector[10] = fifoOut[9][11];
              muxOutConnector[11] = fifoOut[10][11];
              muxOutConnector[12] = fifoOut[11][11];
              muxOutConnector[13] = fifoOut[12][11];
              muxOutConnector[14] = fifoOut[13][11];
              muxOutConnector[15] = fifoOut[14][11];
              muxOutConnector[16] = fifoOut[15][11];
              muxOutConnector[17] = fifoOut[16][11];
              muxOutConnector[18] = fifoOut[17][11];
              muxOutConnector[19] = fifoOut[18][11];
              muxOutConnector[20] = fifoOut[19][11];
              muxOutConnector[21] = fifoOut[20][11];
              muxOutConnector[22] = fifoOut[21][11];
              muxOutConnector[23] = fifoOut[22][11];
              muxOutConnector[24] = fifoOut[23][11];
              muxOutConnector[25] = fifoOut[24][11];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       15: begin
              muxOutConnector[0] = fifoOut[25][12];
              muxOutConnector[1] = fifoOut[0][11];
              muxOutConnector[2] = fifoOut[1][11];
              muxOutConnector[3] = fifoOut[2][11];
              muxOutConnector[4] = fifoOut[3][11];
              muxOutConnector[5] = fifoOut[4][11];
              muxOutConnector[6] = fifoOut[5][11];
              muxOutConnector[7] = fifoOut[6][11];
              muxOutConnector[8] = fifoOut[7][11];
              muxOutConnector[9] = fifoOut[8][11];
              muxOutConnector[10] = fifoOut[9][11];
              muxOutConnector[11] = fifoOut[10][11];
              muxOutConnector[12] = fifoOut[11][11];
              muxOutConnector[13] = fifoOut[12][11];
              muxOutConnector[14] = fifoOut[13][11];
              muxOutConnector[15] = fifoOut[14][11];
              muxOutConnector[16] = fifoOut[15][11];
              muxOutConnector[17] = fifoOut[16][11];
              muxOutConnector[18] = fifoOut[17][11];
              muxOutConnector[19] = fifoOut[18][11];
              muxOutConnector[20] = fifoOut[19][11];
              muxOutConnector[21] = fifoOut[20][11];
              muxOutConnector[22] = fifoOut[21][11];
              muxOutConnector[23] = fifoOut[22][11];
              muxOutConnector[24] = fifoOut[23][11];
              muxOutConnector[25] = fifoOut[24][11];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       16: begin
              muxOutConnector[0] = fifoOut[25][12];
              muxOutConnector[1] = fifoOut[0][11];
              muxOutConnector[2] = fifoOut[1][11];
              muxOutConnector[3] = fifoOut[2][11];
              muxOutConnector[4] = fifoOut[3][11];
              muxOutConnector[5] = fifoOut[4][11];
              muxOutConnector[6] = fifoOut[5][11];
              muxOutConnector[7] = fifoOut[6][11];
              muxOutConnector[8] = fifoOut[7][11];
              muxOutConnector[9] = fifoOut[8][11];
              muxOutConnector[10] = fifoOut[9][11];
              muxOutConnector[11] = fifoOut[10][11];
              muxOutConnector[12] = fifoOut[11][11];
              muxOutConnector[13] = fifoOut[12][11];
              muxOutConnector[14] = fifoOut[13][11];
              muxOutConnector[15] = fifoOut[14][11];
              muxOutConnector[16] = fifoOut[15][11];
              muxOutConnector[17] = fifoOut[16][11];
              muxOutConnector[18] = fifoOut[17][11];
              muxOutConnector[19] = fifoOut[18][11];
              muxOutConnector[20] = fifoOut[19][11];
              muxOutConnector[21] = fifoOut[20][11];
              muxOutConnector[22] = fifoOut[21][11];
              muxOutConnector[23] = fifoOut[22][11];
              muxOutConnector[24] = fifoOut[23][11];
              muxOutConnector[25] = fifoOut[24][11];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       17: begin
              muxOutConnector[0] = fifoOut[25][12];
              muxOutConnector[1] = fifoOut[0][11];
              muxOutConnector[2] = fifoOut[1][11];
              muxOutConnector[3] = fifoOut[2][11];
              muxOutConnector[4] = fifoOut[3][11];
              muxOutConnector[5] = fifoOut[4][11];
              muxOutConnector[6] = fifoOut[5][11];
              muxOutConnector[7] = fifoOut[6][11];
              muxOutConnector[8] = fifoOut[7][11];
              muxOutConnector[9] = fifoOut[8][11];
              muxOutConnector[10] = fifoOut[9][11];
              muxOutConnector[11] = fifoOut[10][11];
              muxOutConnector[12] = fifoOut[11][11];
              muxOutConnector[13] = fifoOut[12][11];
              muxOutConnector[14] = fifoOut[13][11];
              muxOutConnector[15] = fifoOut[14][11];
              muxOutConnector[16] = fifoOut[15][11];
              muxOutConnector[17] = fifoOut[16][11];
              muxOutConnector[18] = fifoOut[17][11];
              muxOutConnector[19] = fifoOut[18][11];
              muxOutConnector[20] = fifoOut[19][11];
              muxOutConnector[21] = fifoOut[20][11];
              muxOutConnector[22] = fifoOut[21][11];
              muxOutConnector[23] = fifoOut[22][11];
              muxOutConnector[24] = fifoOut[23][11];
              muxOutConnector[25] = fifoOut[24][11];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       18: begin
              muxOutConnector[0] = fifoOut[25][12];
              muxOutConnector[1] = fifoOut[0][11];
              muxOutConnector[2] = fifoOut[1][11];
              muxOutConnector[3] = fifoOut[2][11];
              muxOutConnector[4] = fifoOut[3][11];
              muxOutConnector[5] = fifoOut[4][11];
              muxOutConnector[6] = fifoOut[5][11];
              muxOutConnector[7] = fifoOut[6][11];
              muxOutConnector[8] = fifoOut[7][11];
              muxOutConnector[9] = fifoOut[8][11];
              muxOutConnector[10] = fifoOut[9][11];
              muxOutConnector[11] = fifoOut[10][11];
              muxOutConnector[12] = fifoOut[11][11];
              muxOutConnector[13] = fifoOut[12][11];
              muxOutConnector[14] = fifoOut[13][11];
              muxOutConnector[15] = fifoOut[14][11];
              muxOutConnector[16] = fifoOut[15][11];
              muxOutConnector[17] = fifoOut[16][11];
              muxOutConnector[18] = fifoOut[17][11];
              muxOutConnector[19] = fifoOut[18][11];
              muxOutConnector[20] = fifoOut[19][11];
              muxOutConnector[21] = fifoOut[20][11];
              muxOutConnector[22] = fifoOut[21][11];
              muxOutConnector[23] = fifoOut[22][11];
              muxOutConnector[24] = fifoOut[23][11];
              muxOutConnector[25] = fifoOut[24][11];
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = fifoOut[49][9];
              muxOutConnector[44] = fifoOut[50][9];
              muxOutConnector[45] = fifoOut[51][9];
              muxOutConnector[46] = fifoOut[26][8];
              muxOutConnector[47] = fifoOut[27][8];
              muxOutConnector[48] = fifoOut[28][8];
              muxOutConnector[49] = fifoOut[29][8];
              muxOutConnector[50] = fifoOut[30][8];
              muxOutConnector[51] = fifoOut[31][8];
       end
       19: begin
              muxOutConnector[0] = fifoOut[25][12];
              muxOutConnector[1] = fifoOut[0][11];
              muxOutConnector[2] = fifoOut[1][11];
              muxOutConnector[3] = fifoOut[2][11];
              muxOutConnector[4] = fifoOut[3][11];
              muxOutConnector[5] = fifoOut[4][11];
              muxOutConnector[6] = fifoOut[5][11];
              muxOutConnector[7] = fifoOut[6][11];
              muxOutConnector[8] = fifoOut[7][11];
              muxOutConnector[9] = fifoOut[8][11];
              muxOutConnector[10] = fifoOut[9][11];
              muxOutConnector[11] = fifoOut[10][11];
              muxOutConnector[12] = fifoOut[11][11];
              muxOutConnector[13] = fifoOut[12][11];
              muxOutConnector[14] = fifoOut[13][11];
              muxOutConnector[15] = fifoOut[14][11];
              muxOutConnector[16] = fifoOut[15][11];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[32][9];
              muxOutConnector[27] = fifoOut[33][9];
              muxOutConnector[28] = fifoOut[34][9];
              muxOutConnector[29] = fifoOut[35][9];
              muxOutConnector[30] = fifoOut[36][9];
              muxOutConnector[31] = fifoOut[37][9];
              muxOutConnector[32] = fifoOut[38][9];
              muxOutConnector[33] = fifoOut[39][9];
              muxOutConnector[34] = fifoOut[40][9];
              muxOutConnector[35] = fifoOut[41][9];
              muxOutConnector[36] = fifoOut[42][9];
              muxOutConnector[37] = fifoOut[43][9];
              muxOutConnector[38] = fifoOut[44][9];
              muxOutConnector[39] = fifoOut[45][9];
              muxOutConnector[40] = fifoOut[46][9];
              muxOutConnector[41] = fifoOut[47][9];
              muxOutConnector[42] = fifoOut[48][9];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
