`timescale 1ns / 1ps
module LMem1To0_511_circ2_combined_ys_yu_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        rxIn,
        load_input_en,
        iteration_0_indicator,
        feedback_en,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter r_lower = 32;
parameter c = 17;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input load_input_en;
input iteration_0_indicator;
input [ADDRESSWIDTH-1:0]unloadAddress;
input feedback_en;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input [ r_lower * w - 1 : 0 ] rxIn; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
wire [w-1:0]rxInConnector[r_lower-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

generate
    for (k=0;k<r_lower;k=k+1)begin:assign_rx
        assign rxInConnector[k] = rxIn[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            if(feedback_en)begin
                 fifoOut[i][0] <= fifoOut[i][c-1];
            end
            else if(load_input_en)begin
                 if(i < r_lower)begin
                   fifoOut[i][0] = rxInConnector[i];
                 end
                 else begin
                   fifoOut[i][0] = maxVal;
                 end
            end
            else begin
                 fifoOut[i][0] <= ly0InConnector[i];
            end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
       0: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = fifoOut[1][7][w-1];
              unloadMuxOut[31] = fifoOut[2][7][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[3][8][w-1];
              unloadMuxOut[1] = fifoOut[4][8][w-1];
              unloadMuxOut[2] = fifoOut[5][8][w-1];
              unloadMuxOut[3] = fifoOut[6][8][w-1];
              unloadMuxOut[4] = fifoOut[7][8][w-1];
              unloadMuxOut[5] = fifoOut[8][8][w-1];
              unloadMuxOut[6] = fifoOut[9][8][w-1];
              unloadMuxOut[7] = fifoOut[10][8][w-1];
              unloadMuxOut[8] = fifoOut[11][8][w-1];
              unloadMuxOut[9] = fifoOut[12][8][w-1];
              unloadMuxOut[10] = fifoOut[13][8][w-1];
              unloadMuxOut[11] = fifoOut[14][8][w-1];
              unloadMuxOut[12] = fifoOut[15][8][w-1];
              unloadMuxOut[13] = fifoOut[16][8][w-1];
              unloadMuxOut[14] = fifoOut[17][8][w-1];
              unloadMuxOut[15] = fifoOut[18][8][w-1];
              unloadMuxOut[16] = fifoOut[19][8][w-1];
              unloadMuxOut[17] = fifoOut[20][8][w-1];
              unloadMuxOut[18] = fifoOut[21][8][w-1];
              unloadMuxOut[19] = fifoOut[22][8][w-1];
              unloadMuxOut[20] = fifoOut[23][8][w-1];
              unloadMuxOut[21] = fifoOut[24][8][w-1];
              unloadMuxOut[22] = fifoOut[25][8][w-1];
              unloadMuxOut[23] = fifoOut[0][7][w-1];
              unloadMuxOut[24] = fifoOut[1][7][w-1];
              unloadMuxOut[25] = fifoOut[2][7][w-1];
              unloadMuxOut[26] = fifoOut[3][7][w-1];
              unloadMuxOut[27] = fifoOut[4][7][w-1];
              unloadMuxOut[28] = fifoOut[5][7][w-1];
              unloadMuxOut[29] = fifoOut[6][7][w-1];
              unloadMuxOut[30] = fifoOut[7][7][w-1];
              unloadMuxOut[31] = fifoOut[8][7][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[9][8][w-1];
              unloadMuxOut[1] = fifoOut[10][8][w-1];
              unloadMuxOut[2] = fifoOut[11][8][w-1];
              unloadMuxOut[3] = fifoOut[12][8][w-1];
              unloadMuxOut[4] = fifoOut[13][8][w-1];
              unloadMuxOut[5] = fifoOut[14][8][w-1];
              unloadMuxOut[6] = fifoOut[15][8][w-1];
              unloadMuxOut[7] = fifoOut[16][8][w-1];
              unloadMuxOut[8] = fifoOut[17][8][w-1];
              unloadMuxOut[9] = fifoOut[18][8][w-1];
              unloadMuxOut[10] = fifoOut[19][8][w-1];
              unloadMuxOut[11] = fifoOut[20][8][w-1];
              unloadMuxOut[12] = fifoOut[21][8][w-1];
              unloadMuxOut[13] = fifoOut[22][8][w-1];
              unloadMuxOut[14] = fifoOut[23][8][w-1];
              unloadMuxOut[15] = fifoOut[24][8][w-1];
              unloadMuxOut[16] = fifoOut[25][8][w-1];
              unloadMuxOut[17] = fifoOut[0][7][w-1];
              unloadMuxOut[18] = fifoOut[1][7][w-1];
              unloadMuxOut[19] = fifoOut[2][7][w-1];
              unloadMuxOut[20] = fifoOut[3][7][w-1];
              unloadMuxOut[21] = fifoOut[4][7][w-1];
              unloadMuxOut[22] = fifoOut[5][7][w-1];
              unloadMuxOut[23] = fifoOut[6][7][w-1];
              unloadMuxOut[24] = fifoOut[7][7][w-1];
              unloadMuxOut[25] = fifoOut[8][7][w-1];
              unloadMuxOut[26] = fifoOut[9][7][w-1];
              unloadMuxOut[27] = fifoOut[10][7][w-1];
              unloadMuxOut[28] = fifoOut[11][7][w-1];
              unloadMuxOut[29] = fifoOut[12][7][w-1];
              unloadMuxOut[30] = fifoOut[13][7][w-1];
              unloadMuxOut[31] = fifoOut[14][7][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[15][8][w-1];
              unloadMuxOut[1] = fifoOut[16][8][w-1];
              unloadMuxOut[2] = fifoOut[17][8][w-1];
              unloadMuxOut[3] = fifoOut[18][8][w-1];
              unloadMuxOut[4] = fifoOut[19][8][w-1];
              unloadMuxOut[5] = fifoOut[20][8][w-1];
              unloadMuxOut[6] = fifoOut[21][8][w-1];
              unloadMuxOut[7] = fifoOut[22][8][w-1];
              unloadMuxOut[8] = fifoOut[23][8][w-1];
              unloadMuxOut[9] = fifoOut[24][8][w-1];
              unloadMuxOut[10] = fifoOut[25][8][w-1];
              unloadMuxOut[11] = fifoOut[0][7][w-1];
              unloadMuxOut[12] = fifoOut[1][7][w-1];
              unloadMuxOut[13] = fifoOut[2][7][w-1];
              unloadMuxOut[14] = fifoOut[3][7][w-1];
              unloadMuxOut[15] = fifoOut[4][7][w-1];
              unloadMuxOut[16] = fifoOut[5][7][w-1];
              unloadMuxOut[17] = fifoOut[6][7][w-1];
              unloadMuxOut[18] = fifoOut[7][7][w-1];
              unloadMuxOut[19] = fifoOut[8][7][w-1];
              unloadMuxOut[20] = fifoOut[9][7][w-1];
              unloadMuxOut[21] = fifoOut[10][7][w-1];
              unloadMuxOut[22] = fifoOut[11][7][w-1];
              unloadMuxOut[23] = fifoOut[12][7][w-1];
              unloadMuxOut[24] = fifoOut[13][7][w-1];
              unloadMuxOut[25] = fifoOut[14][7][w-1];
              unloadMuxOut[26] = fifoOut[15][7][w-1];
              unloadMuxOut[27] = fifoOut[16][7][w-1];
              unloadMuxOut[28] = fifoOut[17][7][w-1];
              unloadMuxOut[29] = fifoOut[18][7][w-1];
              unloadMuxOut[30] = fifoOut[19][7][w-1];
              unloadMuxOut[31] = fifoOut[20][7][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[21][8][w-1];
              unloadMuxOut[1] = fifoOut[22][8][w-1];
              unloadMuxOut[2] = fifoOut[23][8][w-1];
              unloadMuxOut[3] = fifoOut[24][8][w-1];
              unloadMuxOut[4] = fifoOut[25][8][w-1];
              unloadMuxOut[5] = fifoOut[0][7][w-1];
              unloadMuxOut[6] = fifoOut[1][7][w-1];
              unloadMuxOut[7] = fifoOut[2][7][w-1];
              unloadMuxOut[8] = fifoOut[3][7][w-1];
              unloadMuxOut[9] = fifoOut[4][7][w-1];
              unloadMuxOut[10] = fifoOut[5][7][w-1];
              unloadMuxOut[11] = fifoOut[6][7][w-1];
              unloadMuxOut[12] = fifoOut[7][7][w-1];
              unloadMuxOut[13] = fifoOut[8][7][w-1];
              unloadMuxOut[14] = fifoOut[9][7][w-1];
              unloadMuxOut[15] = fifoOut[10][7][w-1];
              unloadMuxOut[16] = fifoOut[11][7][w-1];
              unloadMuxOut[17] = fifoOut[12][7][w-1];
              unloadMuxOut[18] = fifoOut[13][7][w-1];
              unloadMuxOut[19] = fifoOut[14][7][w-1];
              unloadMuxOut[20] = fifoOut[15][7][w-1];
              unloadMuxOut[21] = fifoOut[16][7][w-1];
              unloadMuxOut[22] = fifoOut[17][7][w-1];
              unloadMuxOut[23] = fifoOut[18][7][w-1];
              unloadMuxOut[24] = fifoOut[19][7][w-1];
              unloadMuxOut[25] = fifoOut[20][7][w-1];
              unloadMuxOut[26] = fifoOut[21][7][w-1];
              unloadMuxOut[27] = fifoOut[22][7][w-1];
              unloadMuxOut[28] = fifoOut[23][7][w-1];
              unloadMuxOut[29] = fifoOut[24][7][w-1];
              unloadMuxOut[30] = fifoOut[25][7][w-1];
              unloadMuxOut[31] = fifoOut[0][6][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[1][7][w-1];
              unloadMuxOut[1] = fifoOut[2][7][w-1];
              unloadMuxOut[2] = fifoOut[3][7][w-1];
              unloadMuxOut[3] = fifoOut[4][7][w-1];
              unloadMuxOut[4] = fifoOut[5][7][w-1];
              unloadMuxOut[5] = fifoOut[6][7][w-1];
              unloadMuxOut[6] = fifoOut[7][7][w-1];
              unloadMuxOut[7] = fifoOut[8][7][w-1];
              unloadMuxOut[8] = fifoOut[9][7][w-1];
              unloadMuxOut[9] = fifoOut[10][7][w-1];
              unloadMuxOut[10] = fifoOut[11][7][w-1];
              unloadMuxOut[11] = fifoOut[12][7][w-1];
              unloadMuxOut[12] = fifoOut[13][7][w-1];
              unloadMuxOut[13] = fifoOut[14][7][w-1];
              unloadMuxOut[14] = fifoOut[15][7][w-1];
              unloadMuxOut[15] = fifoOut[16][7][w-1];
              unloadMuxOut[16] = fifoOut[17][7][w-1];
              unloadMuxOut[17] = fifoOut[18][7][w-1];
              unloadMuxOut[18] = fifoOut[19][7][w-1];
              unloadMuxOut[19] = fifoOut[20][7][w-1];
              unloadMuxOut[20] = fifoOut[21][7][w-1];
              unloadMuxOut[21] = fifoOut[22][7][w-1];
              unloadMuxOut[22] = fifoOut[23][7][w-1];
              unloadMuxOut[23] = fifoOut[24][7][w-1];
              unloadMuxOut[24] = fifoOut[25][7][w-1];
              unloadMuxOut[25] = fifoOut[0][6][w-1];
              unloadMuxOut[26] = fifoOut[1][6][w-1];
              unloadMuxOut[27] = fifoOut[2][6][w-1];
              unloadMuxOut[28] = fifoOut[26][15][w-1];
              unloadMuxOut[29] = fifoOut[27][15][w-1];
              unloadMuxOut[30] = fifoOut[28][15][w-1];
              unloadMuxOut[31] = fifoOut[29][15][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[30][16][w-1];
              unloadMuxOut[1] = fifoOut[31][16][w-1];
              unloadMuxOut[2] = fifoOut[32][16][w-1];
              unloadMuxOut[3] = fifoOut[33][16][w-1];
              unloadMuxOut[4] = fifoOut[34][16][w-1];
              unloadMuxOut[5] = fifoOut[35][16][w-1];
              unloadMuxOut[6] = fifoOut[36][16][w-1];
              unloadMuxOut[7] = fifoOut[37][16][w-1];
              unloadMuxOut[8] = fifoOut[38][16][w-1];
              unloadMuxOut[9] = fifoOut[39][16][w-1];
              unloadMuxOut[10] = fifoOut[40][16][w-1];
              unloadMuxOut[11] = fifoOut[41][16][w-1];
              unloadMuxOut[12] = fifoOut[42][16][w-1];
              unloadMuxOut[13] = fifoOut[43][16][w-1];
              unloadMuxOut[14] = fifoOut[44][16][w-1];
              unloadMuxOut[15] = fifoOut[45][16][w-1];
              unloadMuxOut[16] = fifoOut[46][16][w-1];
              unloadMuxOut[17] = fifoOut[47][16][w-1];
              unloadMuxOut[18] = fifoOut[48][16][w-1];
              unloadMuxOut[19] = fifoOut[49][16][w-1];
              unloadMuxOut[20] = fifoOut[50][16][w-1];
              unloadMuxOut[21] = fifoOut[51][16][w-1];
              unloadMuxOut[22] = fifoOut[26][15][w-1];
              unloadMuxOut[23] = fifoOut[27][15][w-1];
              unloadMuxOut[24] = fifoOut[28][15][w-1];
              unloadMuxOut[25] = fifoOut[29][15][w-1];
              unloadMuxOut[26] = fifoOut[30][15][w-1];
              unloadMuxOut[27] = fifoOut[31][15][w-1];
              unloadMuxOut[28] = fifoOut[32][15][w-1];
              unloadMuxOut[29] = fifoOut[33][15][w-1];
              unloadMuxOut[30] = fifoOut[34][15][w-1];
              unloadMuxOut[31] = fifoOut[35][15][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[36][16][w-1];
              unloadMuxOut[1] = fifoOut[37][16][w-1];
              unloadMuxOut[2] = fifoOut[38][16][w-1];
              unloadMuxOut[3] = fifoOut[39][16][w-1];
              unloadMuxOut[4] = fifoOut[40][16][w-1];
              unloadMuxOut[5] = fifoOut[41][16][w-1];
              unloadMuxOut[6] = fifoOut[42][16][w-1];
              unloadMuxOut[7] = fifoOut[43][16][w-1];
              unloadMuxOut[8] = fifoOut[44][16][w-1];
              unloadMuxOut[9] = fifoOut[45][16][w-1];
              unloadMuxOut[10] = fifoOut[46][16][w-1];
              unloadMuxOut[11] = fifoOut[47][16][w-1];
              unloadMuxOut[12] = fifoOut[48][16][w-1];
              unloadMuxOut[13] = fifoOut[49][16][w-1];
              unloadMuxOut[14] = fifoOut[50][16][w-1];
              unloadMuxOut[15] = fifoOut[51][16][w-1];
              unloadMuxOut[16] = fifoOut[26][15][w-1];
              unloadMuxOut[17] = fifoOut[27][15][w-1];
              unloadMuxOut[18] = fifoOut[28][15][w-1];
              unloadMuxOut[19] = fifoOut[29][15][w-1];
              unloadMuxOut[20] = fifoOut[30][15][w-1];
              unloadMuxOut[21] = fifoOut[31][15][w-1];
              unloadMuxOut[22] = fifoOut[32][15][w-1];
              unloadMuxOut[23] = fifoOut[33][15][w-1];
              unloadMuxOut[24] = fifoOut[34][15][w-1];
              unloadMuxOut[25] = fifoOut[35][15][w-1];
              unloadMuxOut[26] = fifoOut[36][15][w-1];
              unloadMuxOut[27] = fifoOut[37][15][w-1];
              unloadMuxOut[28] = fifoOut[38][15][w-1];
              unloadMuxOut[29] = fifoOut[39][15][w-1];
              unloadMuxOut[30] = fifoOut[40][15][w-1];
              unloadMuxOut[31] = fifoOut[41][15][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[42][16][w-1];
              unloadMuxOut[1] = fifoOut[43][16][w-1];
              unloadMuxOut[2] = fifoOut[44][16][w-1];
              unloadMuxOut[3] = fifoOut[45][16][w-1];
              unloadMuxOut[4] = fifoOut[46][16][w-1];
              unloadMuxOut[5] = fifoOut[47][16][w-1];
              unloadMuxOut[6] = fifoOut[48][16][w-1];
              unloadMuxOut[7] = fifoOut[49][16][w-1];
              unloadMuxOut[8] = fifoOut[50][16][w-1];
              unloadMuxOut[9] = fifoOut[51][16][w-1];
              unloadMuxOut[10] = fifoOut[26][15][w-1];
              unloadMuxOut[11] = fifoOut[27][15][w-1];
              unloadMuxOut[12] = fifoOut[28][15][w-1];
              unloadMuxOut[13] = fifoOut[29][15][w-1];
              unloadMuxOut[14] = fifoOut[30][15][w-1];
              unloadMuxOut[15] = fifoOut[31][15][w-1];
              unloadMuxOut[16] = fifoOut[32][15][w-1];
              unloadMuxOut[17] = fifoOut[33][15][w-1];
              unloadMuxOut[18] = fifoOut[34][15][w-1];
              unloadMuxOut[19] = fifoOut[35][15][w-1];
              unloadMuxOut[20] = fifoOut[36][15][w-1];
              unloadMuxOut[21] = fifoOut[37][15][w-1];
              unloadMuxOut[22] = fifoOut[38][15][w-1];
              unloadMuxOut[23] = fifoOut[39][15][w-1];
              unloadMuxOut[24] = fifoOut[40][15][w-1];
              unloadMuxOut[25] = fifoOut[41][15][w-1];
              unloadMuxOut[26] = fifoOut[42][15][w-1];
              unloadMuxOut[27] = fifoOut[43][15][w-1];
              unloadMuxOut[28] = fifoOut[44][15][w-1];
              unloadMuxOut[29] = fifoOut[45][15][w-1];
              unloadMuxOut[30] = fifoOut[46][15][w-1];
              unloadMuxOut[31] = fifoOut[47][15][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[48][16][w-1];
              unloadMuxOut[1] = fifoOut[49][16][w-1];
              unloadMuxOut[2] = fifoOut[50][16][w-1];
              unloadMuxOut[3] = fifoOut[51][16][w-1];
              unloadMuxOut[4] = fifoOut[26][15][w-1];
              unloadMuxOut[5] = fifoOut[27][15][w-1];
              unloadMuxOut[6] = fifoOut[28][15][w-1];
              unloadMuxOut[7] = fifoOut[29][15][w-1];
              unloadMuxOut[8] = fifoOut[30][15][w-1];
              unloadMuxOut[9] = fifoOut[31][15][w-1];
              unloadMuxOut[10] = fifoOut[32][15][w-1];
              unloadMuxOut[11] = fifoOut[33][15][w-1];
              unloadMuxOut[12] = fifoOut[34][15][w-1];
              unloadMuxOut[13] = fifoOut[35][15][w-1];
              unloadMuxOut[14] = fifoOut[36][15][w-1];
              unloadMuxOut[15] = fifoOut[37][15][w-1];
              unloadMuxOut[16] = fifoOut[38][15][w-1];
              unloadMuxOut[17] = fifoOut[39][15][w-1];
              unloadMuxOut[18] = fifoOut[40][15][w-1];
              unloadMuxOut[19] = fifoOut[41][15][w-1];
              unloadMuxOut[20] = fifoOut[42][15][w-1];
              unloadMuxOut[21] = fifoOut[43][15][w-1];
              unloadMuxOut[22] = fifoOut[44][15][w-1];
              unloadMuxOut[23] = fifoOut[45][15][w-1];
              unloadMuxOut[24] = fifoOut[46][15][w-1];
              unloadMuxOut[25] = fifoOut[47][15][w-1];
              unloadMuxOut[26] = fifoOut[48][15][w-1];
              unloadMuxOut[27] = fifoOut[49][15][w-1];
              unloadMuxOut[28] = fifoOut[50][15][w-1];
              unloadMuxOut[29] = fifoOut[51][15][w-1];
              unloadMuxOut[30] = fifoOut[26][14][w-1];
              unloadMuxOut[31] = fifoOut[27][14][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[28][15][w-1];
              unloadMuxOut[1] = fifoOut[29][15][w-1];
              unloadMuxOut[2] = fifoOut[30][15][w-1];
              unloadMuxOut[3] = fifoOut[31][15][w-1];
              unloadMuxOut[4] = fifoOut[32][15][w-1];
              unloadMuxOut[5] = fifoOut[33][15][w-1];
              unloadMuxOut[6] = fifoOut[34][15][w-1];
              unloadMuxOut[7] = fifoOut[35][15][w-1];
              unloadMuxOut[8] = fifoOut[36][15][w-1];
              unloadMuxOut[9] = fifoOut[37][15][w-1];
              unloadMuxOut[10] = fifoOut[38][15][w-1];
              unloadMuxOut[11] = fifoOut[39][15][w-1];
              unloadMuxOut[12] = fifoOut[40][15][w-1];
              unloadMuxOut[13] = fifoOut[41][15][w-1];
              unloadMuxOut[14] = fifoOut[42][15][w-1];
              unloadMuxOut[15] = fifoOut[43][15][w-1];
              unloadMuxOut[16] = fifoOut[44][15][w-1];
              unloadMuxOut[17] = fifoOut[45][15][w-1];
              unloadMuxOut[18] = fifoOut[46][15][w-1];
              unloadMuxOut[19] = fifoOut[47][15][w-1];
              unloadMuxOut[20] = fifoOut[48][15][w-1];
              unloadMuxOut[21] = fifoOut[49][15][w-1];
              unloadMuxOut[22] = fifoOut[50][15][w-1];
              unloadMuxOut[23] = fifoOut[51][15][w-1];
              unloadMuxOut[24] = fifoOut[26][14][w-1];
              unloadMuxOut[25] = fifoOut[27][14][w-1];
              unloadMuxOut[26] = fifoOut[28][14][w-1];
              unloadMuxOut[27] = fifoOut[29][14][w-1];
              unloadMuxOut[28] = fifoOut[30][14][w-1];
              unloadMuxOut[29] = fifoOut[31][14][w-1];
              unloadMuxOut[30] = fifoOut[32][14][w-1];
              unloadMuxOut[31] = fifoOut[33][14][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[34][15][w-1];
              unloadMuxOut[1] = fifoOut[35][15][w-1];
              unloadMuxOut[2] = fifoOut[36][15][w-1];
              unloadMuxOut[3] = fifoOut[37][15][w-1];
              unloadMuxOut[4] = fifoOut[38][15][w-1];
              unloadMuxOut[5] = fifoOut[39][15][w-1];
              unloadMuxOut[6] = fifoOut[40][15][w-1];
              unloadMuxOut[7] = fifoOut[41][15][w-1];
              unloadMuxOut[8] = fifoOut[42][15][w-1];
              unloadMuxOut[9] = fifoOut[43][15][w-1];
              unloadMuxOut[10] = fifoOut[44][15][w-1];
              unloadMuxOut[11] = fifoOut[45][15][w-1];
              unloadMuxOut[12] = fifoOut[46][15][w-1];
              unloadMuxOut[13] = fifoOut[47][15][w-1];
              unloadMuxOut[14] = fifoOut[48][15][w-1];
              unloadMuxOut[15] = fifoOut[49][15][w-1];
              unloadMuxOut[16] = fifoOut[50][15][w-1];
              unloadMuxOut[17] = fifoOut[51][15][w-1];
              unloadMuxOut[18] = fifoOut[26][14][w-1];
              unloadMuxOut[19] = fifoOut[27][14][w-1];
              unloadMuxOut[20] = fifoOut[28][14][w-1];
              unloadMuxOut[21] = fifoOut[29][14][w-1];
              unloadMuxOut[22] = fifoOut[30][14][w-1];
              unloadMuxOut[23] = fifoOut[31][14][w-1];
              unloadMuxOut[24] = fifoOut[32][14][w-1];
              unloadMuxOut[25] = fifoOut[33][14][w-1];
              unloadMuxOut[26] = fifoOut[34][14][w-1];
              unloadMuxOut[27] = fifoOut[35][14][w-1];
              unloadMuxOut[28] = fifoOut[36][14][w-1];
              unloadMuxOut[29] = fifoOut[37][14][w-1];
              unloadMuxOut[30] = fifoOut[38][14][w-1];
              unloadMuxOut[31] = fifoOut[39][14][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[40][15][w-1];
              unloadMuxOut[1] = fifoOut[41][15][w-1];
              unloadMuxOut[2] = fifoOut[42][15][w-1];
              unloadMuxOut[3] = fifoOut[43][15][w-1];
              unloadMuxOut[4] = fifoOut[44][15][w-1];
              unloadMuxOut[5] = fifoOut[45][15][w-1];
              unloadMuxOut[6] = fifoOut[46][15][w-1];
              unloadMuxOut[7] = fifoOut[47][15][w-1];
              unloadMuxOut[8] = fifoOut[48][15][w-1];
              unloadMuxOut[9] = fifoOut[49][15][w-1];
              unloadMuxOut[10] = fifoOut[50][15][w-1];
              unloadMuxOut[11] = fifoOut[51][15][w-1];
              unloadMuxOut[12] = fifoOut[26][14][w-1];
              unloadMuxOut[13] = fifoOut[27][14][w-1];
              unloadMuxOut[14] = fifoOut[28][14][w-1];
              unloadMuxOut[15] = fifoOut[29][14][w-1];
              unloadMuxOut[16] = fifoOut[30][14][w-1];
              unloadMuxOut[17] = fifoOut[31][14][w-1];
              unloadMuxOut[18] = fifoOut[32][14][w-1];
              unloadMuxOut[19] = fifoOut[33][14][w-1];
              unloadMuxOut[20] = fifoOut[34][14][w-1];
              unloadMuxOut[21] = fifoOut[35][14][w-1];
              unloadMuxOut[22] = fifoOut[36][14][w-1];
              unloadMuxOut[23] = fifoOut[37][14][w-1];
              unloadMuxOut[24] = fifoOut[38][14][w-1];
              unloadMuxOut[25] = fifoOut[39][14][w-1];
              unloadMuxOut[26] = fifoOut[40][14][w-1];
              unloadMuxOut[27] = fifoOut[41][14][w-1];
              unloadMuxOut[28] = fifoOut[42][14][w-1];
              unloadMuxOut[29] = fifoOut[43][14][w-1];
              unloadMuxOut[30] = fifoOut[44][14][w-1];
              unloadMuxOut[31] = fifoOut[45][14][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[46][15][w-1];
              unloadMuxOut[1] = fifoOut[47][15][w-1];
              unloadMuxOut[2] = fifoOut[48][15][w-1];
              unloadMuxOut[3] = fifoOut[49][15][w-1];
              unloadMuxOut[4] = fifoOut[50][15][w-1];
              unloadMuxOut[5] = fifoOut[51][15][w-1];
              unloadMuxOut[6] = fifoOut[26][14][w-1];
              unloadMuxOut[7] = fifoOut[27][14][w-1];
              unloadMuxOut[8] = fifoOut[28][14][w-1];
              unloadMuxOut[9] = fifoOut[29][14][w-1];
              unloadMuxOut[10] = fifoOut[30][14][w-1];
              unloadMuxOut[11] = fifoOut[31][14][w-1];
              unloadMuxOut[12] = fifoOut[32][14][w-1];
              unloadMuxOut[13] = fifoOut[33][14][w-1];
              unloadMuxOut[14] = fifoOut[34][14][w-1];
              unloadMuxOut[15] = fifoOut[35][14][w-1];
              unloadMuxOut[16] = fifoOut[36][14][w-1];
              unloadMuxOut[17] = fifoOut[37][14][w-1];
              unloadMuxOut[18] = fifoOut[38][14][w-1];
              unloadMuxOut[19] = fifoOut[39][14][w-1];
              unloadMuxOut[20] = fifoOut[40][14][w-1];
              unloadMuxOut[21] = fifoOut[41][14][w-1];
              unloadMuxOut[22] = fifoOut[42][14][w-1];
              unloadMuxOut[23] = fifoOut[43][14][w-1];
              unloadMuxOut[24] = fifoOut[44][14][w-1];
              unloadMuxOut[25] = fifoOut[45][14][w-1];
              unloadMuxOut[26] = fifoOut[46][14][w-1];
              unloadMuxOut[27] = fifoOut[47][14][w-1];
              unloadMuxOut[28] = fifoOut[48][14][w-1];
              unloadMuxOut[29] = fifoOut[49][14][w-1];
              unloadMuxOut[30] = fifoOut[50][14][w-1];
              unloadMuxOut[31] = fifoOut[51][14][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[26][14][w-1];
              unloadMuxOut[1] = fifoOut[27][14][w-1];
              unloadMuxOut[2] = fifoOut[28][14][w-1];
              unloadMuxOut[3] = fifoOut[29][14][w-1];
              unloadMuxOut[4] = fifoOut[30][14][w-1];
              unloadMuxOut[5] = fifoOut[31][14][w-1];
              unloadMuxOut[6] = fifoOut[32][14][w-1];
              unloadMuxOut[7] = fifoOut[33][14][w-1];
              unloadMuxOut[8] = fifoOut[34][14][w-1];
              unloadMuxOut[9] = fifoOut[35][14][w-1];
              unloadMuxOut[10] = fifoOut[36][14][w-1];
              unloadMuxOut[11] = fifoOut[37][14][w-1];
              unloadMuxOut[12] = fifoOut[38][14][w-1];
              unloadMuxOut[13] = fifoOut[39][14][w-1];
              unloadMuxOut[14] = fifoOut[40][14][w-1];
              unloadMuxOut[15] = fifoOut[41][14][w-1];
              unloadMuxOut[16] = fifoOut[42][14][w-1];
              unloadMuxOut[17] = fifoOut[3][7][w-1];
              unloadMuxOut[18] = fifoOut[4][7][w-1];
              unloadMuxOut[19] = fifoOut[5][7][w-1];
              unloadMuxOut[20] = fifoOut[6][7][w-1];
              unloadMuxOut[21] = fifoOut[7][7][w-1];
              unloadMuxOut[22] = fifoOut[8][7][w-1];
              unloadMuxOut[23] = fifoOut[9][7][w-1];
              unloadMuxOut[24] = fifoOut[10][7][w-1];
              unloadMuxOut[25] = fifoOut[11][7][w-1];
              unloadMuxOut[26] = fifoOut[12][7][w-1];
              unloadMuxOut[27] = fifoOut[13][7][w-1];
              unloadMuxOut[28] = fifoOut[14][7][w-1];
              unloadMuxOut[29] = fifoOut[15][7][w-1];
              unloadMuxOut[30] = fifoOut[16][7][w-1];
              unloadMuxOut[31] = fifoOut[17][7][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[18][8][w-1];
              unloadMuxOut[1] = fifoOut[19][8][w-1];
              unloadMuxOut[2] = fifoOut[20][8][w-1];
              unloadMuxOut[3] = fifoOut[21][8][w-1];
              unloadMuxOut[4] = fifoOut[22][8][w-1];
              unloadMuxOut[5] = fifoOut[23][8][w-1];
              unloadMuxOut[6] = fifoOut[24][8][w-1];
              unloadMuxOut[7] = fifoOut[25][8][w-1];
              unloadMuxOut[8] = fifoOut[0][7][w-1];
              unloadMuxOut[9] = fifoOut[1][7][w-1];
              unloadMuxOut[10] = fifoOut[2][7][w-1];
              unloadMuxOut[11] = fifoOut[3][7][w-1];
              unloadMuxOut[12] = fifoOut[4][7][w-1];
              unloadMuxOut[13] = fifoOut[5][7][w-1];
              unloadMuxOut[14] = fifoOut[6][7][w-1];
              unloadMuxOut[15] = fifoOut[7][7][w-1];
              unloadMuxOut[16] = fifoOut[8][7][w-1];
              unloadMuxOut[17] = fifoOut[9][7][w-1];
              unloadMuxOut[18] = fifoOut[10][7][w-1];
              unloadMuxOut[19] = fifoOut[11][7][w-1];
              unloadMuxOut[20] = fifoOut[12][7][w-1];
              unloadMuxOut[21] = fifoOut[13][7][w-1];
              unloadMuxOut[22] = fifoOut[14][7][w-1];
              unloadMuxOut[23] = fifoOut[15][7][w-1];
              unloadMuxOut[24] = fifoOut[16][7][w-1];
              unloadMuxOut[25] = fifoOut[17][7][w-1];
              unloadMuxOut[26] = fifoOut[18][7][w-1];
              unloadMuxOut[27] = fifoOut[19][7][w-1];
              unloadMuxOut[28] = fifoOut[20][7][w-1];
              unloadMuxOut[29] = fifoOut[21][7][w-1];
              unloadMuxOut[30] = fifoOut[22][7][w-1];
              unloadMuxOut[31] = fifoOut[23][7][w-1];
       end
       16: begin
              unloadMuxOut[0] = fifoOut[24][8][w-1];
              unloadMuxOut[1] = fifoOut[25][8][w-1];
              unloadMuxOut[2] = fifoOut[0][7][w-1];
              unloadMuxOut[3] = fifoOut[1][7][w-1];
              unloadMuxOut[4] = fifoOut[2][7][w-1];
              unloadMuxOut[5] = fifoOut[3][7][w-1];
              unloadMuxOut[6] = fifoOut[4][7][w-1];
              unloadMuxOut[7] = fifoOut[5][7][w-1];
              unloadMuxOut[8] = fifoOut[6][7][w-1];
              unloadMuxOut[9] = fifoOut[7][7][w-1];
              unloadMuxOut[10] = fifoOut[8][7][w-1];
              unloadMuxOut[11] = fifoOut[9][7][w-1];
              unloadMuxOut[12] = fifoOut[10][7][w-1];
              unloadMuxOut[13] = fifoOut[11][7][w-1];
              unloadMuxOut[14] = fifoOut[12][7][w-1];
              unloadMuxOut[15] = fifoOut[13][7][w-1];
              unloadMuxOut[16] = fifoOut[14][7][w-1];
              unloadMuxOut[17] = fifoOut[15][7][w-1];
              unloadMuxOut[18] = fifoOut[16][7][w-1];
              unloadMuxOut[19] = fifoOut[17][7][w-1];
              unloadMuxOut[20] = fifoOut[18][7][w-1];
              unloadMuxOut[21] = fifoOut[19][7][w-1];
              unloadMuxOut[22] = fifoOut[20][7][w-1];
              unloadMuxOut[23] = fifoOut[21][7][w-1];
              unloadMuxOut[24] = fifoOut[22][7][w-1];
              unloadMuxOut[25] = fifoOut[23][7][w-1];
              unloadMuxOut[26] = fifoOut[24][7][w-1];
              unloadMuxOut[27] = fifoOut[25][7][w-1];
              unloadMuxOut[28] = fifoOut[0][6][w-1];
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0; 
             end
       end
    endcase //unload case end
    case(iteration_0_indicator)
       0: begin
         case(rd_address_case)
         0: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[38][3];
              muxOutConnector[27] = fifoOut[39][3];
              muxOutConnector[28] = fifoOut[40][3];
              muxOutConnector[29] = fifoOut[41][3];
              muxOutConnector[30] = fifoOut[42][3];
              muxOutConnector[31] = fifoOut[43][3];
              muxOutConnector[32] = fifoOut[44][3];
              muxOutConnector[33] = fifoOut[45][3];
              muxOutConnector[34] = fifoOut[46][3];
              muxOutConnector[35] = fifoOut[47][3];
              muxOutConnector[36] = fifoOut[48][3];
              muxOutConnector[37] = fifoOut[49][3];
              muxOutConnector[38] = fifoOut[50][3];
              muxOutConnector[39] = fifoOut[51][3];
              muxOutConnector[40] = fifoOut[26][2];
              muxOutConnector[41] = fifoOut[27][2];
              muxOutConnector[42] = fifoOut[28][2];
              muxOutConnector[43] = fifoOut[29][2];
              muxOutConnector[44] = fifoOut[30][2];
              muxOutConnector[45] = fifoOut[31][2];
              muxOutConnector[46] = fifoOut[32][2];
              muxOutConnector[47] = fifoOut[33][2];
              muxOutConnector[48] = fifoOut[34][2];
              muxOutConnector[49] = fifoOut[35][2];
              muxOutConnector[50] = fifoOut[36][2];
              muxOutConnector[51] = fifoOut[37][2];
         end
         1: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[38][3];
              muxOutConnector[27] = fifoOut[39][3];
              muxOutConnector[28] = fifoOut[40][3];
              muxOutConnector[29] = fifoOut[41][3];
              muxOutConnector[30] = fifoOut[42][3];
              muxOutConnector[31] = fifoOut[43][3];
              muxOutConnector[32] = fifoOut[44][3];
              muxOutConnector[33] = fifoOut[45][3];
              muxOutConnector[34] = fifoOut[46][3];
              muxOutConnector[35] = fifoOut[47][3];
              muxOutConnector[36] = fifoOut[48][3];
              muxOutConnector[37] = fifoOut[49][3];
              muxOutConnector[38] = fifoOut[50][3];
              muxOutConnector[39] = fifoOut[51][3];
              muxOutConnector[40] = fifoOut[26][2];
              muxOutConnector[41] = fifoOut[27][2];
              muxOutConnector[42] = fifoOut[28][2];
              muxOutConnector[43] = fifoOut[29][2];
              muxOutConnector[44] = fifoOut[30][2];
              muxOutConnector[45] = fifoOut[31][2];
              muxOutConnector[46] = fifoOut[32][2];
              muxOutConnector[47] = fifoOut[33][2];
              muxOutConnector[48] = fifoOut[34][2];
              muxOutConnector[49] = fifoOut[35][2];
              muxOutConnector[50] = fifoOut[36][2];
              muxOutConnector[51] = fifoOut[37][2];
         end
         2: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[38][3];
              muxOutConnector[27] = fifoOut[39][3];
              muxOutConnector[28] = fifoOut[40][3];
              muxOutConnector[29] = fifoOut[41][3];
              muxOutConnector[30] = fifoOut[42][3];
              muxOutConnector[31] = fifoOut[43][3];
              muxOutConnector[32] = fifoOut[44][3];
              muxOutConnector[33] = fifoOut[45][3];
              muxOutConnector[34] = fifoOut[46][3];
              muxOutConnector[35] = fifoOut[47][3];
              muxOutConnector[36] = fifoOut[48][3];
              muxOutConnector[37] = fifoOut[49][3];
              muxOutConnector[38] = fifoOut[50][3];
              muxOutConnector[39] = fifoOut[51][3];
              muxOutConnector[40] = fifoOut[26][2];
              muxOutConnector[41] = fifoOut[27][2];
              muxOutConnector[42] = fifoOut[28][2];
              muxOutConnector[43] = fifoOut[29][2];
              muxOutConnector[44] = fifoOut[30][2];
              muxOutConnector[45] = fifoOut[31][2];
              muxOutConnector[46] = fifoOut[32][2];
              muxOutConnector[47] = fifoOut[33][2];
              muxOutConnector[48] = fifoOut[34][2];
              muxOutConnector[49] = fifoOut[35][2];
              muxOutConnector[50] = fifoOut[36][2];
              muxOutConnector[51] = fifoOut[37][2];
         end
         3: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[38][3];
              muxOutConnector[27] = fifoOut[39][3];
              muxOutConnector[28] = fifoOut[0][13];
              muxOutConnector[29] = fifoOut[1][13];
              muxOutConnector[30] = fifoOut[2][13];
              muxOutConnector[31] = fifoOut[3][13];
              muxOutConnector[32] = fifoOut[4][13];
              muxOutConnector[33] = fifoOut[5][13];
              muxOutConnector[34] = fifoOut[6][13];
              muxOutConnector[35] = fifoOut[7][13];
              muxOutConnector[36] = fifoOut[8][13];
              muxOutConnector[37] = fifoOut[9][13];
              muxOutConnector[38] = fifoOut[10][13];
              muxOutConnector[39] = fifoOut[11][13];
              muxOutConnector[40] = fifoOut[12][13];
              muxOutConnector[41] = fifoOut[13][13];
              muxOutConnector[42] = fifoOut[14][13];
              muxOutConnector[43] = fifoOut[15][13];
              muxOutConnector[44] = fifoOut[16][13];
              muxOutConnector[45] = fifoOut[17][13];
              muxOutConnector[46] = fifoOut[18][13];
              muxOutConnector[47] = fifoOut[19][13];
              muxOutConnector[48] = fifoOut[20][13];
              muxOutConnector[49] = fifoOut[21][13];
              muxOutConnector[50] = fifoOut[22][13];
              muxOutConnector[51] = fifoOut[23][13];
         end
         4: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[24][14];
              muxOutConnector[27] = fifoOut[25][14];
              muxOutConnector[28] = fifoOut[0][13];
              muxOutConnector[29] = fifoOut[1][13];
              muxOutConnector[30] = fifoOut[2][13];
              muxOutConnector[31] = fifoOut[3][13];
              muxOutConnector[32] = fifoOut[4][13];
              muxOutConnector[33] = fifoOut[5][13];
              muxOutConnector[34] = fifoOut[6][13];
              muxOutConnector[35] = fifoOut[7][13];
              muxOutConnector[36] = fifoOut[8][13];
              muxOutConnector[37] = fifoOut[9][13];
              muxOutConnector[38] = fifoOut[10][13];
              muxOutConnector[39] = fifoOut[11][13];
              muxOutConnector[40] = fifoOut[12][13];
              muxOutConnector[41] = fifoOut[13][13];
              muxOutConnector[42] = fifoOut[14][13];
              muxOutConnector[43] = fifoOut[15][13];
              muxOutConnector[44] = fifoOut[16][13];
              muxOutConnector[45] = fifoOut[17][13];
              muxOutConnector[46] = fifoOut[18][13];
              muxOutConnector[47] = fifoOut[19][13];
              muxOutConnector[48] = fifoOut[20][13];
              muxOutConnector[49] = fifoOut[21][13];
              muxOutConnector[50] = fifoOut[22][13];
              muxOutConnector[51] = fifoOut[23][13];
         end
         5: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[24][14];
              muxOutConnector[27] = fifoOut[25][14];
              muxOutConnector[28] = fifoOut[0][13];
              muxOutConnector[29] = fifoOut[1][13];
              muxOutConnector[30] = fifoOut[2][13];
              muxOutConnector[31] = fifoOut[3][13];
              muxOutConnector[32] = fifoOut[4][13];
              muxOutConnector[33] = fifoOut[5][13];
              muxOutConnector[34] = fifoOut[6][13];
              muxOutConnector[35] = fifoOut[7][13];
              muxOutConnector[36] = fifoOut[8][13];
              muxOutConnector[37] = fifoOut[9][13];
              muxOutConnector[38] = fifoOut[10][13];
              muxOutConnector[39] = fifoOut[11][13];
              muxOutConnector[40] = fifoOut[12][13];
              muxOutConnector[41] = fifoOut[13][13];
              muxOutConnector[42] = fifoOut[14][13];
              muxOutConnector[43] = fifoOut[15][13];
              muxOutConnector[44] = fifoOut[16][13];
              muxOutConnector[45] = fifoOut[17][13];
              muxOutConnector[46] = fifoOut[18][13];
              muxOutConnector[47] = fifoOut[19][13];
              muxOutConnector[48] = fifoOut[20][13];
              muxOutConnector[49] = fifoOut[21][13];
              muxOutConnector[50] = fifoOut[22][13];
              muxOutConnector[51] = fifoOut[23][13];
         end
         6: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[26][16];
              muxOutConnector[3] = fifoOut[27][16];
              muxOutConnector[4] = fifoOut[28][16];
              muxOutConnector[5] = fifoOut[29][16];
              muxOutConnector[6] = fifoOut[30][16];
              muxOutConnector[7] = fifoOut[31][16];
              muxOutConnector[8] = fifoOut[32][16];
              muxOutConnector[9] = fifoOut[33][16];
              muxOutConnector[10] = fifoOut[34][16];
              muxOutConnector[11] = fifoOut[35][16];
              muxOutConnector[12] = fifoOut[36][16];
              muxOutConnector[13] = fifoOut[37][16];
              muxOutConnector[14] = fifoOut[38][16];
              muxOutConnector[15] = fifoOut[39][16];
              muxOutConnector[16] = fifoOut[40][16];
              muxOutConnector[17] = fifoOut[41][16];
              muxOutConnector[18] = fifoOut[42][16];
              muxOutConnector[19] = fifoOut[43][16];
              muxOutConnector[20] = fifoOut[44][16];
              muxOutConnector[21] = fifoOut[45][16];
              muxOutConnector[22] = fifoOut[46][16];
              muxOutConnector[23] = fifoOut[47][16];
              muxOutConnector[24] = fifoOut[48][16];
              muxOutConnector[25] = fifoOut[49][16];
              muxOutConnector[26] = fifoOut[24][14];
              muxOutConnector[27] = fifoOut[25][14];
              muxOutConnector[28] = fifoOut[0][13];
              muxOutConnector[29] = fifoOut[1][13];
              muxOutConnector[30] = fifoOut[2][13];
              muxOutConnector[31] = fifoOut[3][13];
              muxOutConnector[32] = fifoOut[4][13];
              muxOutConnector[33] = fifoOut[5][13];
              muxOutConnector[34] = fifoOut[6][13];
              muxOutConnector[35] = fifoOut[7][13];
              muxOutConnector[36] = fifoOut[8][13];
              muxOutConnector[37] = fifoOut[9][13];
              muxOutConnector[38] = fifoOut[10][13];
              muxOutConnector[39] = fifoOut[11][13];
              muxOutConnector[40] = fifoOut[12][13];
              muxOutConnector[41] = fifoOut[13][13];
              muxOutConnector[42] = fifoOut[14][13];
              muxOutConnector[43] = fifoOut[15][13];
              muxOutConnector[44] = fifoOut[16][13];
              muxOutConnector[45] = fifoOut[17][13];
              muxOutConnector[46] = fifoOut[18][13];
              muxOutConnector[47] = fifoOut[19][13];
              muxOutConnector[48] = fifoOut[20][13];
              muxOutConnector[49] = fifoOut[21][13];
              muxOutConnector[50] = fifoOut[22][13];
              muxOutConnector[51] = fifoOut[23][13];
         end
         7: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[26][16];
              muxOutConnector[3] = fifoOut[27][16];
              muxOutConnector[4] = fifoOut[28][16];
              muxOutConnector[5] = fifoOut[29][16];
              muxOutConnector[6] = fifoOut[30][16];
              muxOutConnector[7] = fifoOut[31][16];
              muxOutConnector[8] = fifoOut[32][16];
              muxOutConnector[9] = fifoOut[33][16];
              muxOutConnector[10] = fifoOut[34][16];
              muxOutConnector[11] = fifoOut[35][16];
              muxOutConnector[12] = fifoOut[36][16];
              muxOutConnector[13] = fifoOut[37][16];
              muxOutConnector[14] = fifoOut[38][16];
              muxOutConnector[15] = fifoOut[39][16];
              muxOutConnector[16] = fifoOut[40][16];
              muxOutConnector[17] = fifoOut[41][16];
              muxOutConnector[18] = fifoOut[42][16];
              muxOutConnector[19] = fifoOut[43][16];
              muxOutConnector[20] = fifoOut[44][16];
              muxOutConnector[21] = fifoOut[45][16];
              muxOutConnector[22] = fifoOut[46][16];
              muxOutConnector[23] = fifoOut[47][16];
              muxOutConnector[24] = fifoOut[48][16];
              muxOutConnector[25] = fifoOut[49][16];
              muxOutConnector[26] = fifoOut[24][14];
              muxOutConnector[27] = fifoOut[25][14];
              muxOutConnector[28] = fifoOut[0][13];
              muxOutConnector[29] = fifoOut[1][13];
              muxOutConnector[30] = fifoOut[2][13];
              muxOutConnector[31] = fifoOut[3][13];
              muxOutConnector[32] = fifoOut[4][13];
              muxOutConnector[33] = fifoOut[5][13];
              muxOutConnector[34] = fifoOut[6][13];
              muxOutConnector[35] = fifoOut[7][13];
              muxOutConnector[36] = fifoOut[8][13];
              muxOutConnector[37] = fifoOut[9][13];
              muxOutConnector[38] = fifoOut[10][13];
              muxOutConnector[39] = fifoOut[11][13];
              muxOutConnector[40] = fifoOut[12][13];
              muxOutConnector[41] = fifoOut[13][13];
              muxOutConnector[42] = fifoOut[14][13];
              muxOutConnector[43] = fifoOut[15][13];
              muxOutConnector[44] = fifoOut[16][13];
              muxOutConnector[45] = fifoOut[17][13];
              muxOutConnector[46] = fifoOut[18][13];
              muxOutConnector[47] = fifoOut[19][13];
              muxOutConnector[48] = fifoOut[20][13];
              muxOutConnector[49] = fifoOut[21][13];
              muxOutConnector[50] = fifoOut[22][13];
              muxOutConnector[51] = fifoOut[23][13];
         end
         8: begin
              muxOutConnector[0] = fifoOut[50][0];
              muxOutConnector[1] = fifoOut[51][0];
              muxOutConnector[2] = fifoOut[26][16];
              muxOutConnector[3] = fifoOut[27][16];
              muxOutConnector[4] = fifoOut[28][16];
              muxOutConnector[5] = fifoOut[29][16];
              muxOutConnector[6] = fifoOut[30][16];
              muxOutConnector[7] = fifoOut[31][16];
              muxOutConnector[8] = fifoOut[32][16];
              muxOutConnector[9] = fifoOut[33][16];
              muxOutConnector[10] = fifoOut[34][16];
              muxOutConnector[11] = fifoOut[35][16];
              muxOutConnector[12] = fifoOut[36][16];
              muxOutConnector[13] = fifoOut[37][16];
              muxOutConnector[14] = fifoOut[38][16];
              muxOutConnector[15] = fifoOut[39][16];
              muxOutConnector[16] = fifoOut[40][16];
              muxOutConnector[17] = fifoOut[41][16];
              muxOutConnector[18] = fifoOut[42][16];
              muxOutConnector[19] = fifoOut[43][16];
              muxOutConnector[20] = fifoOut[44][16];
              muxOutConnector[21] = fifoOut[45][16];
              muxOutConnector[22] = fifoOut[46][16];
              muxOutConnector[23] = fifoOut[47][16];
              muxOutConnector[24] = fifoOut[48][16];
              muxOutConnector[25] = fifoOut[49][16];
              muxOutConnector[26] = fifoOut[24][14];
              muxOutConnector[27] = fifoOut[25][14];
              muxOutConnector[28] = fifoOut[0][13];
              muxOutConnector[29] = fifoOut[1][13];
              muxOutConnector[30] = fifoOut[2][13];
              muxOutConnector[31] = fifoOut[3][13];
              muxOutConnector[32] = fifoOut[4][13];
              muxOutConnector[33] = fifoOut[5][13];
              muxOutConnector[34] = fifoOut[6][13];
              muxOutConnector[35] = fifoOut[7][13];
              muxOutConnector[36] = fifoOut[8][13];
              muxOutConnector[37] = fifoOut[9][13];
              muxOutConnector[38] = fifoOut[10][13];
              muxOutConnector[39] = fifoOut[11][13];
              muxOutConnector[40] = fifoOut[12][13];
              muxOutConnector[41] = fifoOut[13][13];
              muxOutConnector[42] = fifoOut[14][13];
              muxOutConnector[43] = fifoOut[15][13];
              muxOutConnector[44] = fifoOut[16][13];
              muxOutConnector[45] = fifoOut[17][13];
              muxOutConnector[46] = fifoOut[18][13];
              muxOutConnector[47] = fifoOut[19][13];
              muxOutConnector[48] = fifoOut[20][13];
              muxOutConnector[49] = fifoOut[21][13];
              muxOutConnector[50] = fifoOut[22][13];
              muxOutConnector[51] = fifoOut[23][13];
         end
         9: begin
              muxOutConnector[0] = fifoOut[50][0];
              muxOutConnector[1] = fifoOut[51][0];
              muxOutConnector[2] = fifoOut[26][16];
              muxOutConnector[3] = fifoOut[27][16];
              muxOutConnector[4] = fifoOut[28][16];
              muxOutConnector[5] = fifoOut[29][16];
              muxOutConnector[6] = fifoOut[30][16];
              muxOutConnector[7] = fifoOut[31][16];
              muxOutConnector[8] = fifoOut[32][16];
              muxOutConnector[9] = fifoOut[33][16];
              muxOutConnector[10] = fifoOut[34][16];
              muxOutConnector[11] = fifoOut[35][16];
              muxOutConnector[12] = fifoOut[36][16];
              muxOutConnector[13] = fifoOut[37][16];
              muxOutConnector[14] = fifoOut[38][16];
              muxOutConnector[15] = fifoOut[39][16];
              muxOutConnector[16] = fifoOut[40][16];
              muxOutConnector[17] = fifoOut[41][16];
              muxOutConnector[18] = fifoOut[42][16];
              muxOutConnector[19] = fifoOut[43][16];
              muxOutConnector[20] = fifoOut[44][16];
              muxOutConnector[21] = fifoOut[45][16];
              muxOutConnector[22] = fifoOut[46][16];
              muxOutConnector[23] = fifoOut[47][16];
              muxOutConnector[24] = fifoOut[48][16];
              muxOutConnector[25] = fifoOut[49][16];
              muxOutConnector[26] = fifoOut[24][14];
              muxOutConnector[27] = fifoOut[25][14];
              muxOutConnector[28] = fifoOut[0][13];
              muxOutConnector[29] = fifoOut[1][13];
              muxOutConnector[30] = fifoOut[2][13];
              muxOutConnector[31] = fifoOut[3][13];
              muxOutConnector[32] = fifoOut[4][13];
              muxOutConnector[33] = fifoOut[5][13];
              muxOutConnector[34] = fifoOut[6][13];
              muxOutConnector[35] = fifoOut[7][13];
              muxOutConnector[36] = fifoOut[8][13];
              muxOutConnector[37] = fifoOut[9][13];
              muxOutConnector[38] = fifoOut[10][13];
              muxOutConnector[39] = fifoOut[11][13];
              muxOutConnector[40] = fifoOut[12][13];
              muxOutConnector[41] = fifoOut[13][13];
              muxOutConnector[42] = fifoOut[14][13];
              muxOutConnector[43] = fifoOut[15][13];
              muxOutConnector[44] = fifoOut[16][13];
              muxOutConnector[45] = fifoOut[17][13];
              muxOutConnector[46] = fifoOut[18][13];
              muxOutConnector[47] = fifoOut[19][13];
              muxOutConnector[48] = fifoOut[20][13];
              muxOutConnector[49] = fifoOut[21][13];
              muxOutConnector[50] = fifoOut[22][13];
              muxOutConnector[51] = fifoOut[23][13];
         end
         10: begin
              muxOutConnector[0] = fifoOut[50][0];
              muxOutConnector[1] = fifoOut[51][0];
              muxOutConnector[2] = fifoOut[26][16];
              muxOutConnector[3] = fifoOut[27][16];
              muxOutConnector[4] = fifoOut[28][16];
              muxOutConnector[5] = fifoOut[29][16];
              muxOutConnector[6] = fifoOut[30][16];
              muxOutConnector[7] = fifoOut[31][16];
              muxOutConnector[8] = fifoOut[32][16];
              muxOutConnector[9] = fifoOut[33][16];
              muxOutConnector[10] = fifoOut[34][16];
              muxOutConnector[11] = fifoOut[35][16];
              muxOutConnector[12] = fifoOut[36][16];
              muxOutConnector[13] = fifoOut[37][16];
              muxOutConnector[14] = fifoOut[38][16];
              muxOutConnector[15] = fifoOut[39][16];
              muxOutConnector[16] = fifoOut[40][16];
              muxOutConnector[17] = fifoOut[41][16];
              muxOutConnector[18] = fifoOut[42][16];
              muxOutConnector[19] = fifoOut[43][16];
              muxOutConnector[20] = fifoOut[44][16];
              muxOutConnector[21] = fifoOut[45][16];
              muxOutConnector[22] = fifoOut[46][16];
              muxOutConnector[23] = fifoOut[47][16];
              muxOutConnector[24] = fifoOut[48][16];
              muxOutConnector[25] = fifoOut[49][16];
              muxOutConnector[26] = fifoOut[24][14];
              muxOutConnector[27] = fifoOut[25][14];
              muxOutConnector[28] = fifoOut[0][13];
              muxOutConnector[29] = fifoOut[1][13];
              muxOutConnector[30] = fifoOut[2][13];
              muxOutConnector[31] = fifoOut[3][13];
              muxOutConnector[32] = fifoOut[4][13];
              muxOutConnector[33] = fifoOut[5][13];
              muxOutConnector[34] = fifoOut[6][13];
              muxOutConnector[35] = fifoOut[7][13];
              muxOutConnector[36] = fifoOut[8][13];
              muxOutConnector[37] = fifoOut[9][13];
              muxOutConnector[38] = fifoOut[10][13];
              muxOutConnector[39] = fifoOut[11][13];
              muxOutConnector[40] = fifoOut[12][13];
              muxOutConnector[41] = fifoOut[13][13];
              muxOutConnector[42] = fifoOut[14][13];
              muxOutConnector[43] = fifoOut[15][13];
              muxOutConnector[44] = fifoOut[16][13];
              muxOutConnector[45] = fifoOut[17][13];
              muxOutConnector[46] = fifoOut[18][13];
              muxOutConnector[47] = fifoOut[19][13];
              muxOutConnector[48] = fifoOut[20][13];
              muxOutConnector[49] = fifoOut[21][13];
              muxOutConnector[50] = fifoOut[22][13];
              muxOutConnector[51] = fifoOut[23][13];
         end
         11: begin
              muxOutConnector[0] = fifoOut[50][0];
              muxOutConnector[1] = fifoOut[51][0];
              muxOutConnector[2] = fifoOut[26][16];
              muxOutConnector[3] = fifoOut[27][16];
              muxOutConnector[4] = fifoOut[28][16];
              muxOutConnector[5] = fifoOut[29][16];
              muxOutConnector[6] = fifoOut[30][16];
              muxOutConnector[7] = fifoOut[31][16];
              muxOutConnector[8] = fifoOut[32][16];
              muxOutConnector[9] = fifoOut[33][16];
              muxOutConnector[10] = fifoOut[34][16];
              muxOutConnector[11] = fifoOut[35][16];
              muxOutConnector[12] = fifoOut[36][16];
              muxOutConnector[13] = fifoOut[37][16];
              muxOutConnector[14] = fifoOut[38][16];
              muxOutConnector[15] = fifoOut[39][16];
              muxOutConnector[16] = fifoOut[40][16];
              muxOutConnector[17] = fifoOut[41][16];
              muxOutConnector[18] = fifoOut[42][16];
              muxOutConnector[19] = fifoOut[43][16];
              muxOutConnector[20] = fifoOut[44][16];
              muxOutConnector[21] = fifoOut[45][16];
              muxOutConnector[22] = fifoOut[46][16];
              muxOutConnector[23] = fifoOut[47][16];
              muxOutConnector[24] = fifoOut[48][16];
              muxOutConnector[25] = fifoOut[49][16];
              muxOutConnector[26] = fifoOut[24][14];
              muxOutConnector[27] = fifoOut[25][14];
              muxOutConnector[28] = fifoOut[0][13];
              muxOutConnector[29] = fifoOut[1][13];
              muxOutConnector[30] = fifoOut[2][13];
              muxOutConnector[31] = fifoOut[3][13];
              muxOutConnector[32] = fifoOut[4][13];
              muxOutConnector[33] = fifoOut[5][13];
              muxOutConnector[34] = fifoOut[6][13];
              muxOutConnector[35] = fifoOut[7][13];
              muxOutConnector[36] = fifoOut[8][13];
              muxOutConnector[37] = fifoOut[9][13];
              muxOutConnector[38] = fifoOut[10][13];
              muxOutConnector[39] = fifoOut[11][13];
              muxOutConnector[40] = fifoOut[12][13];
              muxOutConnector[41] = fifoOut[13][13];
              muxOutConnector[42] = fifoOut[14][13];
              muxOutConnector[43] = fifoOut[15][13];
              muxOutConnector[44] = fifoOut[16][13];
              muxOutConnector[45] = fifoOut[17][13];
              muxOutConnector[46] = fifoOut[18][13];
              muxOutConnector[47] = fifoOut[19][13];
              muxOutConnector[48] = fifoOut[20][13];
              muxOutConnector[49] = fifoOut[21][13];
              muxOutConnector[50] = fifoOut[22][13];
              muxOutConnector[51] = fifoOut[23][13];
         end
         12: begin
              muxOutConnector[0] = fifoOut[50][0];
              muxOutConnector[1] = fifoOut[51][0];
              muxOutConnector[2] = fifoOut[26][16];
              muxOutConnector[3] = fifoOut[27][16];
              muxOutConnector[4] = fifoOut[28][16];
              muxOutConnector[5] = fifoOut[29][16];
              muxOutConnector[6] = fifoOut[30][16];
              muxOutConnector[7] = fifoOut[31][16];
              muxOutConnector[8] = fifoOut[32][16];
              muxOutConnector[9] = fifoOut[33][16];
              muxOutConnector[10] = fifoOut[34][16];
              muxOutConnector[11] = fifoOut[35][16];
              muxOutConnector[12] = fifoOut[36][16];
              muxOutConnector[13] = fifoOut[37][16];
              muxOutConnector[14] = fifoOut[38][16];
              muxOutConnector[15] = fifoOut[39][16];
              muxOutConnector[16] = fifoOut[40][16];
              muxOutConnector[17] = fifoOut[41][16];
              muxOutConnector[18] = fifoOut[42][16];
              muxOutConnector[19] = fifoOut[43][16];
              muxOutConnector[20] = fifoOut[44][16];
              muxOutConnector[21] = fifoOut[45][16];
              muxOutConnector[22] = fifoOut[46][16];
              muxOutConnector[23] = fifoOut[47][16];
              muxOutConnector[24] = fifoOut[48][16];
              muxOutConnector[25] = fifoOut[49][16];
              muxOutConnector[26] = fifoOut[24][14];
              muxOutConnector[27] = fifoOut[25][14];
              muxOutConnector[28] = fifoOut[0][13];
              muxOutConnector[29] = fifoOut[1][13];
              muxOutConnector[30] = fifoOut[2][13];
              muxOutConnector[31] = fifoOut[3][13];
              muxOutConnector[32] = fifoOut[4][13];
              muxOutConnector[33] = fifoOut[5][13];
              muxOutConnector[34] = fifoOut[6][13];
              muxOutConnector[35] = fifoOut[7][13];
              muxOutConnector[36] = fifoOut[8][13];
              muxOutConnector[37] = fifoOut[9][13];
              muxOutConnector[38] = fifoOut[10][13];
              muxOutConnector[39] = fifoOut[11][13];
              muxOutConnector[40] = fifoOut[12][13];
              muxOutConnector[41] = fifoOut[13][13];
              muxOutConnector[42] = fifoOut[14][13];
              muxOutConnector[43] = fifoOut[15][13];
              muxOutConnector[44] = fifoOut[16][13];
              muxOutConnector[45] = fifoOut[17][13];
              muxOutConnector[46] = fifoOut[18][13];
              muxOutConnector[47] = fifoOut[19][13];
              muxOutConnector[48] = fifoOut[20][13];
              muxOutConnector[49] = fifoOut[21][13];
              muxOutConnector[50] = fifoOut[22][13];
              muxOutConnector[51] = fifoOut[23][13];
         end
         13: begin
              muxOutConnector[0] = fifoOut[50][0];
              muxOutConnector[1] = fifoOut[51][0];
              muxOutConnector[2] = fifoOut[26][16];
              muxOutConnector[3] = fifoOut[27][16];
              muxOutConnector[4] = fifoOut[28][16];
              muxOutConnector[5] = fifoOut[29][16];
              muxOutConnector[6] = fifoOut[30][16];
              muxOutConnector[7] = fifoOut[31][16];
              muxOutConnector[8] = fifoOut[32][16];
              muxOutConnector[9] = fifoOut[33][16];
              muxOutConnector[10] = fifoOut[34][16];
              muxOutConnector[11] = fifoOut[35][16];
              muxOutConnector[12] = fifoOut[36][16];
              muxOutConnector[13] = fifoOut[37][16];
              muxOutConnector[14] = fifoOut[38][16];
              muxOutConnector[15] = fifoOut[39][16];
              muxOutConnector[16] = fifoOut[40][16];
              muxOutConnector[17] = fifoOut[41][16];
              muxOutConnector[18] = fifoOut[42][16];
              muxOutConnector[19] = fifoOut[43][16];
              muxOutConnector[20] = fifoOut[44][16];
              muxOutConnector[21] = fifoOut[45][16];
              muxOutConnector[22] = fifoOut[46][16];
              muxOutConnector[23] = fifoOut[47][16];
              muxOutConnector[24] = fifoOut[48][16];
              muxOutConnector[25] = fifoOut[49][16];
              muxOutConnector[26] = fifoOut[24][14];
              muxOutConnector[27] = fifoOut[25][14];
              muxOutConnector[28] = fifoOut[0][13];
              muxOutConnector[29] = fifoOut[1][13];
              muxOutConnector[30] = fifoOut[2][13];
              muxOutConnector[31] = fifoOut[3][13];
              muxOutConnector[32] = fifoOut[4][13];
              muxOutConnector[33] = fifoOut[5][13];
              muxOutConnector[34] = fifoOut[6][13];
              muxOutConnector[35] = fifoOut[7][13];
              muxOutConnector[36] = fifoOut[8][13];
              muxOutConnector[37] = fifoOut[9][13];
              muxOutConnector[38] = fifoOut[10][13];
              muxOutConnector[39] = fifoOut[11][13];
              muxOutConnector[40] = fifoOut[12][13];
              muxOutConnector[41] = fifoOut[13][13];
              muxOutConnector[42] = fifoOut[14][13];
              muxOutConnector[43] = fifoOut[15][13];
              muxOutConnector[44] = fifoOut[16][13];
              muxOutConnector[45] = fifoOut[40][5];
              muxOutConnector[46] = fifoOut[41][5];
              muxOutConnector[47] = fifoOut[42][5];
              muxOutConnector[48] = fifoOut[43][5];
              muxOutConnector[49] = fifoOut[44][5];
              muxOutConnector[50] = fifoOut[45][5];
              muxOutConnector[51] = fifoOut[46][5];
         end
         14: begin
              muxOutConnector[0] = fifoOut[50][0];
              muxOutConnector[1] = fifoOut[51][0];
              muxOutConnector[2] = fifoOut[26][16];
              muxOutConnector[3] = fifoOut[27][16];
              muxOutConnector[4] = fifoOut[28][16];
              muxOutConnector[5] = fifoOut[29][16];
              muxOutConnector[6] = fifoOut[30][16];
              muxOutConnector[7] = fifoOut[31][16];
              muxOutConnector[8] = fifoOut[32][16];
              muxOutConnector[9] = fifoOut[33][16];
              muxOutConnector[10] = fifoOut[34][16];
              muxOutConnector[11] = fifoOut[35][16];
              muxOutConnector[12] = fifoOut[36][16];
              muxOutConnector[13] = fifoOut[37][16];
              muxOutConnector[14] = fifoOut[38][16];
              muxOutConnector[15] = fifoOut[39][16];
              muxOutConnector[16] = fifoOut[40][16];
              muxOutConnector[17] = fifoOut[41][16];
              muxOutConnector[18] = fifoOut[42][16];
              muxOutConnector[19] = fifoOut[43][16];
              muxOutConnector[20] = fifoOut[44][16];
              muxOutConnector[21] = fifoOut[45][16];
              muxOutConnector[22] = fifoOut[46][16];
              muxOutConnector[23] = fifoOut[47][16];
              muxOutConnector[24] = fifoOut[48][16];
              muxOutConnector[25] = fifoOut[49][16];
              muxOutConnector[26] = fifoOut[47][6];
              muxOutConnector[27] = fifoOut[48][6];
              muxOutConnector[28] = fifoOut[49][6];
              muxOutConnector[29] = fifoOut[50][6];
              muxOutConnector[30] = fifoOut[51][6];
              muxOutConnector[31] = fifoOut[26][5];
              muxOutConnector[32] = fifoOut[27][5];
              muxOutConnector[33] = fifoOut[28][5];
              muxOutConnector[34] = fifoOut[29][5];
              muxOutConnector[35] = fifoOut[30][5];
              muxOutConnector[36] = fifoOut[31][5];
              muxOutConnector[37] = fifoOut[32][5];
              muxOutConnector[38] = fifoOut[33][5];
              muxOutConnector[39] = fifoOut[34][5];
              muxOutConnector[40] = fifoOut[35][5];
              muxOutConnector[41] = fifoOut[36][5];
              muxOutConnector[42] = fifoOut[37][5];
              muxOutConnector[43] = fifoOut[38][5];
              muxOutConnector[44] = fifoOut[39][5];
              muxOutConnector[45] = fifoOut[40][5];
              muxOutConnector[46] = fifoOut[41][5];
              muxOutConnector[47] = fifoOut[42][5];
              muxOutConnector[48] = fifoOut[43][5];
              muxOutConnector[49] = fifoOut[44][5];
              muxOutConnector[50] = fifoOut[45][5];
              muxOutConnector[51] = fifoOut[46][5];
         end
         15: begin
              muxOutConnector[0] = fifoOut[50][0];
              muxOutConnector[1] = fifoOut[51][0];
              muxOutConnector[2] = fifoOut[26][16];
              muxOutConnector[3] = fifoOut[27][16];
              muxOutConnector[4] = fifoOut[28][16];
              muxOutConnector[5] = fifoOut[29][16];
              muxOutConnector[6] = fifoOut[30][16];
              muxOutConnector[7] = fifoOut[31][16];
              muxOutConnector[8] = fifoOut[32][16];
              muxOutConnector[9] = fifoOut[33][16];
              muxOutConnector[10] = fifoOut[34][16];
              muxOutConnector[11] = fifoOut[35][16];
              muxOutConnector[12] = fifoOut[36][16];
              muxOutConnector[13] = fifoOut[37][16];
              muxOutConnector[14] = fifoOut[38][16];
              muxOutConnector[15] = fifoOut[39][16];
              muxOutConnector[16] = fifoOut[40][16];
              muxOutConnector[17] = fifoOut[41][16];
              muxOutConnector[18] = fifoOut[42][16];
              muxOutConnector[19] = fifoOut[43][16];
              muxOutConnector[20] = fifoOut[44][16];
              muxOutConnector[21] = fifoOut[45][16];
              muxOutConnector[22] = fifoOut[46][16];
              muxOutConnector[23] = fifoOut[47][16];
              muxOutConnector[24] = fifoOut[48][16];
              muxOutConnector[25] = fifoOut[49][16];
              muxOutConnector[26] = fifoOut[47][6];
              muxOutConnector[27] = fifoOut[48][6];
              muxOutConnector[28] = fifoOut[49][6];
              muxOutConnector[29] = fifoOut[50][6];
              muxOutConnector[30] = fifoOut[51][6];
              muxOutConnector[31] = fifoOut[26][5];
              muxOutConnector[32] = fifoOut[27][5];
              muxOutConnector[33] = fifoOut[28][5];
              muxOutConnector[34] = fifoOut[29][5];
              muxOutConnector[35] = fifoOut[30][5];
              muxOutConnector[36] = fifoOut[31][5];
              muxOutConnector[37] = fifoOut[32][5];
              muxOutConnector[38] = fifoOut[33][5];
              muxOutConnector[39] = fifoOut[34][5];
              muxOutConnector[40] = fifoOut[35][5];
              muxOutConnector[41] = fifoOut[36][5];
              muxOutConnector[42] = fifoOut[37][5];
              muxOutConnector[43] = fifoOut[38][5];
              muxOutConnector[44] = fifoOut[39][5];
              muxOutConnector[45] = fifoOut[40][5];
              muxOutConnector[46] = fifoOut[41][5];
              muxOutConnector[47] = fifoOut[42][5];
              muxOutConnector[48] = fifoOut[43][5];
              muxOutConnector[49] = fifoOut[44][5];
              muxOutConnector[50] = fifoOut[45][5];
              muxOutConnector[51] = fifoOut[46][5];
         end
         16: begin
              muxOutConnector[0] = fifoOut[50][0];
              muxOutConnector[1] = fifoOut[51][0];
              muxOutConnector[2] = fifoOut[26][16];
              muxOutConnector[3] = fifoOut[27][16];
              muxOutConnector[4] = fifoOut[28][16];
              muxOutConnector[5] = fifoOut[29][16];
              muxOutConnector[6] = fifoOut[30][16];
              muxOutConnector[7] = fifoOut[31][16];
              muxOutConnector[8] = fifoOut[32][16];
              muxOutConnector[9] = fifoOut[33][16];
              muxOutConnector[10] = fifoOut[34][16];
              muxOutConnector[11] = fifoOut[35][16];
              muxOutConnector[12] = fifoOut[36][16];
              muxOutConnector[13] = fifoOut[37][16];
              muxOutConnector[14] = fifoOut[38][16];
              muxOutConnector[15] = fifoOut[39][16];
              muxOutConnector[16] = fifoOut[40][16];
              muxOutConnector[17] = fifoOut[41][16];
              muxOutConnector[18] = fifoOut[42][16];
              muxOutConnector[19] = fifoOut[3][9];
              muxOutConnector[20] = fifoOut[4][9];
              muxOutConnector[21] = fifoOut[5][9];
              muxOutConnector[22] = fifoOut[6][9];
              muxOutConnector[23] = fifoOut[7][9];
              muxOutConnector[24] = fifoOut[8][9];
              muxOutConnector[25] = fifoOut[9][9];
              muxOutConnector[26] = fifoOut[47][6];
              muxOutConnector[27] = fifoOut[48][6];
              muxOutConnector[28] = fifoOut[49][6];
              muxOutConnector[29] = fifoOut[50][6];
              muxOutConnector[30] = fifoOut[51][6];
              muxOutConnector[31] = fifoOut[26][5];
              muxOutConnector[32] = fifoOut[27][5];
              muxOutConnector[33] = fifoOut[28][5];
              muxOutConnector[34] = fifoOut[29][5];
              muxOutConnector[35] = fifoOut[30][5];
              muxOutConnector[36] = fifoOut[31][5];
              muxOutConnector[37] = fifoOut[32][5];
              muxOutConnector[38] = fifoOut[33][5];
              muxOutConnector[39] = fifoOut[34][5];
              muxOutConnector[40] = fifoOut[35][5];
              muxOutConnector[41] = fifoOut[36][5];
              muxOutConnector[42] = fifoOut[37][5];
              muxOutConnector[43] = fifoOut[38][5];
              muxOutConnector[44] = fifoOut[39][5];
              muxOutConnector[45] = fifoOut[40][5];
              muxOutConnector[46] = fifoOut[41][5];
              muxOutConnector[47] = fifoOut[42][5];
              muxOutConnector[48] = fifoOut[43][5];
              muxOutConnector[49] = fifoOut[44][5];
              muxOutConnector[50] = fifoOut[45][5];
              muxOutConnector[51] = fifoOut[46][5];
         end
         17: begin
              muxOutConnector[0] = fifoOut[10][10];
              muxOutConnector[1] = fifoOut[11][10];
              muxOutConnector[2] = fifoOut[12][10];
              muxOutConnector[3] = fifoOut[13][10];
              muxOutConnector[4] = fifoOut[14][10];
              muxOutConnector[5] = fifoOut[15][10];
              muxOutConnector[6] = fifoOut[16][10];
              muxOutConnector[7] = fifoOut[17][10];
              muxOutConnector[8] = fifoOut[18][10];
              muxOutConnector[9] = fifoOut[19][10];
              muxOutConnector[10] = fifoOut[20][10];
              muxOutConnector[11] = fifoOut[21][10];
              muxOutConnector[12] = fifoOut[22][10];
              muxOutConnector[13] = fifoOut[23][10];
              muxOutConnector[14] = fifoOut[24][10];
              muxOutConnector[15] = fifoOut[25][10];
              muxOutConnector[16] = fifoOut[0][9];
              muxOutConnector[17] = fifoOut[1][9];
              muxOutConnector[18] = fifoOut[2][9];
              muxOutConnector[19] = fifoOut[3][9];
              muxOutConnector[20] = fifoOut[4][9];
              muxOutConnector[21] = fifoOut[5][9];
              muxOutConnector[22] = fifoOut[6][9];
              muxOutConnector[23] = fifoOut[7][9];
              muxOutConnector[24] = fifoOut[8][9];
              muxOutConnector[25] = fifoOut[9][9];
              muxOutConnector[26] = fifoOut[47][6];
              muxOutConnector[27] = fifoOut[48][6];
              muxOutConnector[28] = fifoOut[49][6];
              muxOutConnector[29] = fifoOut[50][6];
              muxOutConnector[30] = fifoOut[51][6];
              muxOutConnector[31] = fifoOut[26][5];
              muxOutConnector[32] = fifoOut[27][5];
              muxOutConnector[33] = fifoOut[28][5];
              muxOutConnector[34] = fifoOut[29][5];
              muxOutConnector[35] = fifoOut[30][5];
              muxOutConnector[36] = fifoOut[31][5];
              muxOutConnector[37] = fifoOut[32][5];
              muxOutConnector[38] = fifoOut[33][5];
              muxOutConnector[39] = fifoOut[34][5];
              muxOutConnector[40] = fifoOut[35][5];
              muxOutConnector[41] = fifoOut[36][5];
              muxOutConnector[42] = fifoOut[37][5];
              muxOutConnector[43] = fifoOut[38][5];
              muxOutConnector[44] = fifoOut[39][5];
              muxOutConnector[45] = fifoOut[40][5];
              muxOutConnector[46] = fifoOut[41][5];
              muxOutConnector[47] = fifoOut[42][5];
              muxOutConnector[48] = fifoOut[43][5];
              muxOutConnector[49] = fifoOut[44][5];
              muxOutConnector[50] = fifoOut[45][5];
              muxOutConnector[51] = fifoOut[46][5];
         end
         18: begin
              muxOutConnector[0] = fifoOut[10][10];
              muxOutConnector[1] = fifoOut[11][10];
              muxOutConnector[2] = fifoOut[12][10];
              muxOutConnector[3] = fifoOut[13][10];
              muxOutConnector[4] = fifoOut[14][10];
              muxOutConnector[5] = fifoOut[15][10];
              muxOutConnector[6] = fifoOut[16][10];
              muxOutConnector[7] = fifoOut[17][10];
              muxOutConnector[8] = fifoOut[18][10];
              muxOutConnector[9] = fifoOut[19][10];
              muxOutConnector[10] = fifoOut[20][10];
              muxOutConnector[11] = fifoOut[21][10];
              muxOutConnector[12] = fifoOut[22][10];
              muxOutConnector[13] = fifoOut[23][10];
              muxOutConnector[14] = fifoOut[24][10];
              muxOutConnector[15] = fifoOut[25][10];
              muxOutConnector[16] = fifoOut[0][9];
              muxOutConnector[17] = fifoOut[1][9];
              muxOutConnector[18] = fifoOut[2][9];
              muxOutConnector[19] = fifoOut[3][9];
              muxOutConnector[20] = fifoOut[4][9];
              muxOutConnector[21] = fifoOut[5][9];
              muxOutConnector[22] = fifoOut[6][9];
              muxOutConnector[23] = fifoOut[7][9];
              muxOutConnector[24] = fifoOut[8][9];
              muxOutConnector[25] = fifoOut[9][9];
              muxOutConnector[26] = fifoOut[47][6];
              muxOutConnector[27] = fifoOut[48][6];
              muxOutConnector[28] = fifoOut[49][6];
              muxOutConnector[29] = fifoOut[50][6];
              muxOutConnector[30] = fifoOut[51][6];
              muxOutConnector[31] = fifoOut[26][5];
              muxOutConnector[32] = fifoOut[27][5];
              muxOutConnector[33] = fifoOut[28][5];
              muxOutConnector[34] = fifoOut[29][5];
              muxOutConnector[35] = fifoOut[30][5];
              muxOutConnector[36] = fifoOut[31][5];
              muxOutConnector[37] = fifoOut[32][5];
              muxOutConnector[38] = fifoOut[33][5];
              muxOutConnector[39] = fifoOut[34][5];
              muxOutConnector[40] = fifoOut[35][5];
              muxOutConnector[41] = fifoOut[36][5];
              muxOutConnector[42] = fifoOut[37][5];
              muxOutConnector[43] = fifoOut[38][5];
              muxOutConnector[44] = fifoOut[39][5];
              muxOutConnector[45] = fifoOut[40][5];
              muxOutConnector[46] = fifoOut[41][5];
              muxOutConnector[47] = fifoOut[42][5];
              muxOutConnector[48] = fifoOut[43][5];
              muxOutConnector[49] = fifoOut[44][5];
              muxOutConnector[50] = fifoOut[45][5];
              muxOutConnector[51] = fifoOut[46][5];
         end
         19: begin
              muxOutConnector[0] = fifoOut[10][10];
              muxOutConnector[1] = fifoOut[11][10];
              muxOutConnector[2] = fifoOut[12][10];
              muxOutConnector[3] = fifoOut[13][10];
              muxOutConnector[4] = fifoOut[14][10];
              muxOutConnector[5] = fifoOut[15][10];
              muxOutConnector[6] = fifoOut[16][10];
              muxOutConnector[7] = fifoOut[17][10];
              muxOutConnector[8] = fifoOut[18][10];
              muxOutConnector[9] = fifoOut[19][10];
              muxOutConnector[10] = fifoOut[20][10];
              muxOutConnector[11] = fifoOut[21][10];
              muxOutConnector[12] = fifoOut[22][10];
              muxOutConnector[13] = fifoOut[23][10];
              muxOutConnector[14] = fifoOut[24][10];
              muxOutConnector[15] = fifoOut[25][10];
              muxOutConnector[16] = fifoOut[0][9];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[47][6];
              muxOutConnector[27] = fifoOut[48][6];
              muxOutConnector[28] = fifoOut[49][6];
              muxOutConnector[29] = fifoOut[50][6];
              muxOutConnector[30] = fifoOut[51][6];
              muxOutConnector[31] = fifoOut[26][5];
              muxOutConnector[32] = fifoOut[27][5];
              muxOutConnector[33] = fifoOut[28][5];
              muxOutConnector[34] = fifoOut[29][5];
              muxOutConnector[35] = fifoOut[30][5];
              muxOutConnector[36] = fifoOut[31][5];
              muxOutConnector[37] = fifoOut[32][5];
              muxOutConnector[38] = fifoOut[33][5];
              muxOutConnector[39] = fifoOut[34][5];
              muxOutConnector[40] = fifoOut[35][5];
              muxOutConnector[41] = fifoOut[36][5];
              muxOutConnector[42] = fifoOut[37][5];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
         end
         default: begin
               for(i=0;i<muxOutSymbols;i=i+1)begin
                muxOutConnector[i] = 0;
              end
         end
//hgjhgbuiguigbigbgbgbui
         endcase
    end
endcase
             end
        endmodule