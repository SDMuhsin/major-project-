`timescale 1ns / 1ps

// Scripted using writeselector_ipintf2_script.m
// based on load symbol pattern table rxregtablemod

// rxregtablemod[row,col] is Nbx17 table, Nb=16 for near earth
// wr_address value= col-1 
// wr_en_vec[idx] and wr_address[idx], idx=circulant subunit mem number = row-1

module writeselector_inputintf(wr_en_vec,wr_address_vec,cyclecount,wr_en);
parameter ADDRESSWIDTH = 5;
parameter Nb = 16;//16*511=8176 codeword

parameter CYCLECOUNTWIDTH = 9;//maxcycles=(8160+64)/32)=257, width=ceil(log2(257))=9

output reg[Nb-1:0] wr_en_vec;
output [(Nb*ADDRESSWIDTH)-1:0] wr_address_vec;
input[(CYCLECOUNTWIDTH)-1:0] cyclecount;
input wr_en;

reg[(ADDRESSWIDTH)-1:0] wr_address[Nb-1:0];
genvar i;
generate
    for (i=0;i<Nb;i=i+1)begin:nb_loop
        assign wr_address_vec[ ((i+1)*ADDRESSWIDTH)-1:i*ADDRESSWIDTH]=wr_address[i];
    end
endgenerate

always@(*) begin
  case(cyclecount)
   1: begin
//row=1, col=1, rxregtablemod(row,col)=-1;
         wr_en_vec[0]=1;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   2: begin
//row=1, col=2, rxregtablemod(row,col)=19;
         wr_en_vec[0]=1;
         wr_address[0]=1;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   3: begin
//row=1, col=3, rxregtablemod(row,col)=51;
         wr_en_vec[0]=1;
         wr_address[0]=2;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   4: begin
//row=1, col=4, rxregtablemod(row,col)=83;
         wr_en_vec[0]=1;
         wr_address[0]=3;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   5: begin
//row=1, col=5, rxregtablemod(row,col)=115;
         wr_en_vec[0]=1;
         wr_address[0]=4;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   6: begin
//row=1, col=6, rxregtablemod(row,col)=147;
         wr_en_vec[0]=1;
         wr_address[0]=5;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   7: begin
//row=1, col=7, rxregtablemod(row,col)=179;
         wr_en_vec[0]=1;
         wr_address[0]=6;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   8: begin
//row=1, col=8, rxregtablemod(row,col)=211;
         wr_en_vec[0]=1;
         wr_address[0]=7;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   9: begin
//row=1, col=9, rxregtablemod(row,col)=243;
         wr_en_vec[0]=1;
         wr_address[0]=8;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   10: begin
//row=1, col=10, rxregtablemod(row,col)=275;
         wr_en_vec[0]=1;
         wr_address[0]=9;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   11: begin
//row=1, col=11, rxregtablemod(row,col)=307;
         wr_en_vec[0]=1;
         wr_address[0]=10;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   12: begin
//row=1, col=12, rxregtablemod(row,col)=339;
         wr_en_vec[0]=1;
         wr_address[0]=11;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   13: begin
//row=1, col=13, rxregtablemod(row,col)=371;
         wr_en_vec[0]=1;
         wr_address[0]=12;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   14: begin
//row=1, col=14, rxregtablemod(row,col)=403;
         wr_en_vec[0]=1;
         wr_address[0]=13;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   15: begin
//row=1, col=15, rxregtablemod(row,col)=435;
         wr_en_vec[0]=1;
         wr_address[0]=14;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   16: begin
//row=1, col=16, rxregtablemod(row,col)=467;
         wr_en_vec[0]=1;
         wr_address[0]=15;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   17: begin
//row=2, col=1, rxregtablemod(row,col)=499;
         wr_en_vec[1]=1;
         wr_address[1]=0;
//row=1, col=17, rxregtablemod(i,17)=499;
         wr_en_vec[0]=1;
         wr_address[0]=16;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   18: begin
//row=2, col=2, rxregtablemod(row,col)=531;
         wr_en_vec[1]=1;
         wr_address[1]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   19: begin
//row=2, col=3, rxregtablemod(row,col)=563;
         wr_en_vec[1]=1;
         wr_address[1]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   20: begin
//row=2, col=4, rxregtablemod(row,col)=595;
         wr_en_vec[1]=1;
         wr_address[1]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   21: begin
//row=2, col=5, rxregtablemod(row,col)=627;
         wr_en_vec[1]=1;
         wr_address[1]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   22: begin
//row=2, col=6, rxregtablemod(row,col)=659;
         wr_en_vec[1]=1;
         wr_address[1]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   23: begin
//row=2, col=7, rxregtablemod(row,col)=691;
         wr_en_vec[1]=1;
         wr_address[1]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   24: begin
//row=2, col=8, rxregtablemod(row,col)=723;
         wr_en_vec[1]=1;
         wr_address[1]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   25: begin
//row=2, col=9, rxregtablemod(row,col)=755;
         wr_en_vec[1]=1;
         wr_address[1]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   26: begin
//row=2, col=10, rxregtablemod(row,col)=787;
         wr_en_vec[1]=1;
         wr_address[1]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   27: begin
//row=2, col=11, rxregtablemod(row,col)=819;
         wr_en_vec[1]=1;
         wr_address[1]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   28: begin
//row=2, col=12, rxregtablemod(row,col)=851;
         wr_en_vec[1]=1;
         wr_address[1]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   29: begin
//row=2, col=13, rxregtablemod(row,col)=883;
         wr_en_vec[1]=1;
         wr_address[1]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   30: begin
//row=2, col=14, rxregtablemod(row,col)=915;
         wr_en_vec[1]=1;
         wr_address[1]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   31: begin
//row=2, col=15, rxregtablemod(row,col)=947;
         wr_en_vec[1]=1;
         wr_address[1]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   32: begin
//row=2, col=16, rxregtablemod(row,col)=979;
         wr_en_vec[1]=1;
         wr_address[1]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   33: begin
//row=3, col=1, rxregtablemod(row,col)=1011;
         wr_en_vec[2]=1;
         wr_address[2]=0;
//row=2, col=17, rxregtablemod(i,17)=1011;
         wr_en_vec[1]=1;
         wr_address[1]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   34: begin
//row=3, col=2, rxregtablemod(row,col)=1043;
         wr_en_vec[2]=1;
         wr_address[2]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   35: begin
//row=3, col=3, rxregtablemod(row,col)=1075;
         wr_en_vec[2]=1;
         wr_address[2]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   36: begin
//row=3, col=4, rxregtablemod(row,col)=1107;
         wr_en_vec[2]=1;
         wr_address[2]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   37: begin
//row=3, col=5, rxregtablemod(row,col)=1139;
         wr_en_vec[2]=1;
         wr_address[2]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   38: begin
//row=3, col=6, rxregtablemod(row,col)=1171;
         wr_en_vec[2]=1;
         wr_address[2]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   39: begin
//row=3, col=7, rxregtablemod(row,col)=1203;
         wr_en_vec[2]=1;
         wr_address[2]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   40: begin
//row=3, col=8, rxregtablemod(row,col)=1235;
         wr_en_vec[2]=1;
         wr_address[2]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   41: begin
//row=3, col=9, rxregtablemod(row,col)=1267;
         wr_en_vec[2]=1;
         wr_address[2]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   42: begin
//row=3, col=10, rxregtablemod(row,col)=1299;
         wr_en_vec[2]=1;
         wr_address[2]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   43: begin
//row=3, col=11, rxregtablemod(row,col)=1331;
         wr_en_vec[2]=1;
         wr_address[2]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   44: begin
//row=3, col=12, rxregtablemod(row,col)=1363;
         wr_en_vec[2]=1;
         wr_address[2]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   45: begin
//row=3, col=13, rxregtablemod(row,col)=1395;
         wr_en_vec[2]=1;
         wr_address[2]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   46: begin
//row=3, col=14, rxregtablemod(row,col)=1427;
         wr_en_vec[2]=1;
         wr_address[2]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   47: begin
//row=3, col=15, rxregtablemod(row,col)=1459;
         wr_en_vec[2]=1;
         wr_address[2]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   48: begin
//row=3, col=16, rxregtablemod(row,col)=1491;
         wr_en_vec[2]=1;
         wr_address[2]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   49: begin
//row=4, col=1, rxregtablemod(row,col)=1523;
         wr_en_vec[3]=1;
         wr_address[3]=0;
//row=3, col=17, rxregtablemod(i,17)=1523;
         wr_en_vec[2]=1;
         wr_address[2]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   50: begin
//row=4, col=2, rxregtablemod(row,col)=1555;
         wr_en_vec[3]=1;
         wr_address[3]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   51: begin
//row=4, col=3, rxregtablemod(row,col)=1587;
         wr_en_vec[3]=1;
         wr_address[3]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   52: begin
//row=4, col=4, rxregtablemod(row,col)=1619;
         wr_en_vec[3]=1;
         wr_address[3]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   53: begin
//row=4, col=5, rxregtablemod(row,col)=1651;
         wr_en_vec[3]=1;
         wr_address[3]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   54: begin
//row=4, col=6, rxregtablemod(row,col)=1683;
         wr_en_vec[3]=1;
         wr_address[3]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   55: begin
//row=4, col=7, rxregtablemod(row,col)=1715;
         wr_en_vec[3]=1;
         wr_address[3]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   56: begin
//row=4, col=8, rxregtablemod(row,col)=1747;
         wr_en_vec[3]=1;
         wr_address[3]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   57: begin
//row=4, col=9, rxregtablemod(row,col)=1779;
         wr_en_vec[3]=1;
         wr_address[3]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   58: begin
//row=4, col=10, rxregtablemod(row,col)=1811;
         wr_en_vec[3]=1;
         wr_address[3]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   59: begin
//row=4, col=11, rxregtablemod(row,col)=1843;
         wr_en_vec[3]=1;
         wr_address[3]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   60: begin
//row=4, col=12, rxregtablemod(row,col)=1875;
         wr_en_vec[3]=1;
         wr_address[3]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   61: begin
//row=4, col=13, rxregtablemod(row,col)=1907;
         wr_en_vec[3]=1;
         wr_address[3]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   62: begin
//row=4, col=14, rxregtablemod(row,col)=1939;
         wr_en_vec[3]=1;
         wr_address[3]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   63: begin
//row=4, col=15, rxregtablemod(row,col)=1971;
         wr_en_vec[3]=1;
         wr_address[3]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   64: begin
//row=4, col=16, rxregtablemod(row,col)=2003;
         wr_en_vec[3]=1;
         wr_address[3]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   65: begin
//row=5, col=1, rxregtablemod(row,col)=2035;
         wr_en_vec[4]=1;
         wr_address[4]=0;
//row=4, col=17, rxregtablemod(i,17)=2035;
         wr_en_vec[3]=1;
         wr_address[3]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   66: begin
//row=5, col=2, rxregtablemod(row,col)=2067;
         wr_en_vec[4]=1;
         wr_address[4]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   67: begin
//row=5, col=3, rxregtablemod(row,col)=2099;
         wr_en_vec[4]=1;
         wr_address[4]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   68: begin
//row=5, col=4, rxregtablemod(row,col)=2131;
         wr_en_vec[4]=1;
         wr_address[4]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   69: begin
//row=5, col=5, rxregtablemod(row,col)=2163;
         wr_en_vec[4]=1;
         wr_address[4]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   70: begin
//row=5, col=6, rxregtablemod(row,col)=2195;
         wr_en_vec[4]=1;
         wr_address[4]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   71: begin
//row=5, col=7, rxregtablemod(row,col)=2227;
         wr_en_vec[4]=1;
         wr_address[4]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   72: begin
//row=5, col=8, rxregtablemod(row,col)=2259;
         wr_en_vec[4]=1;
         wr_address[4]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   73: begin
//row=5, col=9, rxregtablemod(row,col)=2291;
         wr_en_vec[4]=1;
         wr_address[4]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   74: begin
//row=5, col=10, rxregtablemod(row,col)=2323;
         wr_en_vec[4]=1;
         wr_address[4]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   75: begin
//row=5, col=11, rxregtablemod(row,col)=2355;
         wr_en_vec[4]=1;
         wr_address[4]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   76: begin
//row=5, col=12, rxregtablemod(row,col)=2387;
         wr_en_vec[4]=1;
         wr_address[4]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   77: begin
//row=5, col=13, rxregtablemod(row,col)=2419;
         wr_en_vec[4]=1;
         wr_address[4]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   78: begin
//row=5, col=14, rxregtablemod(row,col)=2451;
         wr_en_vec[4]=1;
         wr_address[4]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   79: begin
//row=5, col=15, rxregtablemod(row,col)=2483;
         wr_en_vec[4]=1;
         wr_address[4]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   80: begin
//row=5, col=16, rxregtablemod(row,col)=2515;
         wr_en_vec[4]=1;
         wr_address[4]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   81: begin
//row=6, col=1, rxregtablemod(row,col)=2547;
         wr_en_vec[5]=1;
         wr_address[5]=0;
//row=5, col=17, rxregtablemod(i,17)=2547;
         wr_en_vec[4]=1;
         wr_address[4]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   82: begin
//row=6, col=2, rxregtablemod(row,col)=2579;
         wr_en_vec[5]=1;
         wr_address[5]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   83: begin
//row=6, col=3, rxregtablemod(row,col)=2611;
         wr_en_vec[5]=1;
         wr_address[5]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   84: begin
//row=6, col=4, rxregtablemod(row,col)=2643;
         wr_en_vec[5]=1;
         wr_address[5]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   85: begin
//row=6, col=5, rxregtablemod(row,col)=2675;
         wr_en_vec[5]=1;
         wr_address[5]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   86: begin
//row=6, col=6, rxregtablemod(row,col)=2707;
         wr_en_vec[5]=1;
         wr_address[5]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   87: begin
//row=6, col=7, rxregtablemod(row,col)=2739;
         wr_en_vec[5]=1;
         wr_address[5]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   88: begin
//row=6, col=8, rxregtablemod(row,col)=2771;
         wr_en_vec[5]=1;
         wr_address[5]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   89: begin
//row=6, col=9, rxregtablemod(row,col)=2803;
         wr_en_vec[5]=1;
         wr_address[5]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   90: begin
//row=6, col=10, rxregtablemod(row,col)=2835;
         wr_en_vec[5]=1;
         wr_address[5]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   91: begin
//row=6, col=11, rxregtablemod(row,col)=2867;
         wr_en_vec[5]=1;
         wr_address[5]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   92: begin
//row=6, col=12, rxregtablemod(row,col)=2899;
         wr_en_vec[5]=1;
         wr_address[5]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   93: begin
//row=6, col=13, rxregtablemod(row,col)=2931;
         wr_en_vec[5]=1;
         wr_address[5]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   94: begin
//row=6, col=14, rxregtablemod(row,col)=2963;
         wr_en_vec[5]=1;
         wr_address[5]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   95: begin
//row=6, col=15, rxregtablemod(row,col)=2995;
         wr_en_vec[5]=1;
         wr_address[5]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   96: begin
//row=6, col=16, rxregtablemod(row,col)=3027;
         wr_en_vec[5]=1;
         wr_address[5]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   97: begin
//row=7, col=1, rxregtablemod(row,col)=3059;
         wr_en_vec[6]=1;
         wr_address[6]=0;
//row=6, col=17, rxregtablemod(i,17)=3059;
         wr_en_vec[5]=1;
         wr_address[5]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   98: begin
//row=7, col=2, rxregtablemod(row,col)=3091;
         wr_en_vec[6]=1;
         wr_address[6]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   99: begin
//row=7, col=3, rxregtablemod(row,col)=3123;
         wr_en_vec[6]=1;
         wr_address[6]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   100: begin
//row=7, col=4, rxregtablemod(row,col)=3155;
         wr_en_vec[6]=1;
         wr_address[6]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   101: begin
//row=7, col=5, rxregtablemod(row,col)=3187;
         wr_en_vec[6]=1;
         wr_address[6]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   102: begin
//row=7, col=6, rxregtablemod(row,col)=3219;
         wr_en_vec[6]=1;
         wr_address[6]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   103: begin
//row=7, col=7, rxregtablemod(row,col)=3251;
         wr_en_vec[6]=1;
         wr_address[6]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   104: begin
//row=7, col=8, rxregtablemod(row,col)=3283;
         wr_en_vec[6]=1;
         wr_address[6]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   105: begin
//row=7, col=9, rxregtablemod(row,col)=3315;
         wr_en_vec[6]=1;
         wr_address[6]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   106: begin
//row=7, col=10, rxregtablemod(row,col)=3347;
         wr_en_vec[6]=1;
         wr_address[6]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   107: begin
//row=7, col=11, rxregtablemod(row,col)=3379;
         wr_en_vec[6]=1;
         wr_address[6]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   108: begin
//row=7, col=12, rxregtablemod(row,col)=3411;
         wr_en_vec[6]=1;
         wr_address[6]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   109: begin
//row=7, col=13, rxregtablemod(row,col)=3443;
         wr_en_vec[6]=1;
         wr_address[6]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   110: begin
//row=7, col=14, rxregtablemod(row,col)=3475;
         wr_en_vec[6]=1;
         wr_address[6]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   111: begin
//row=7, col=15, rxregtablemod(row,col)=3507;
         wr_en_vec[6]=1;
         wr_address[6]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   112: begin
//row=7, col=16, rxregtablemod(row,col)=3539;
         wr_en_vec[6]=1;
         wr_address[6]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   113: begin
//row=8, col=1, rxregtablemod(row,col)=3571;
         wr_en_vec[7]=1;
         wr_address[7]=0;
//row=7, col=17, rxregtablemod(i,17)=3571;
         wr_en_vec[6]=1;
         wr_address[6]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   114: begin
//row=8, col=2, rxregtablemod(row,col)=3603;
         wr_en_vec[7]=1;
         wr_address[7]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   115: begin
//row=8, col=3, rxregtablemod(row,col)=3635;
         wr_en_vec[7]=1;
         wr_address[7]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   116: begin
//row=8, col=4, rxregtablemod(row,col)=3667;
         wr_en_vec[7]=1;
         wr_address[7]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   117: begin
//row=8, col=5, rxregtablemod(row,col)=3699;
         wr_en_vec[7]=1;
         wr_address[7]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   118: begin
//row=8, col=6, rxregtablemod(row,col)=3731;
         wr_en_vec[7]=1;
         wr_address[7]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   119: begin
//row=8, col=7, rxregtablemod(row,col)=3763;
         wr_en_vec[7]=1;
         wr_address[7]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   120: begin
//row=8, col=8, rxregtablemod(row,col)=3795;
         wr_en_vec[7]=1;
         wr_address[7]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   121: begin
//row=8, col=9, rxregtablemod(row,col)=3827;
         wr_en_vec[7]=1;
         wr_address[7]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   122: begin
//row=8, col=10, rxregtablemod(row,col)=3859;
         wr_en_vec[7]=1;
         wr_address[7]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   123: begin
//row=8, col=11, rxregtablemod(row,col)=3891;
         wr_en_vec[7]=1;
         wr_address[7]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   124: begin
//row=8, col=12, rxregtablemod(row,col)=3923;
         wr_en_vec[7]=1;
         wr_address[7]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   125: begin
//row=8, col=13, rxregtablemod(row,col)=3955;
         wr_en_vec[7]=1;
         wr_address[7]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   126: begin
//row=8, col=14, rxregtablemod(row,col)=3987;
         wr_en_vec[7]=1;
         wr_address[7]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   127: begin
//row=8, col=15, rxregtablemod(row,col)=4019;
         wr_en_vec[7]=1;
         wr_address[7]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   128: begin
//row=8, col=16, rxregtablemod(row,col)=4051;
         wr_en_vec[7]=1;
         wr_address[7]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   129: begin
//row=9, col=1, rxregtablemod(row,col)=4083;
         wr_en_vec[8]=1;
         wr_address[8]=0;
//row=8, col=17, rxregtablemod(i,17)=4083;
         wr_en_vec[7]=1;
         wr_address[7]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   130: begin
//row=9, col=2, rxregtablemod(row,col)=4115;
         wr_en_vec[8]=1;
         wr_address[8]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   131: begin
//row=9, col=3, rxregtablemod(row,col)=4147;
         wr_en_vec[8]=1;
         wr_address[8]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   132: begin
//row=9, col=4, rxregtablemod(row,col)=4179;
         wr_en_vec[8]=1;
         wr_address[8]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   133: begin
//row=9, col=5, rxregtablemod(row,col)=4211;
         wr_en_vec[8]=1;
         wr_address[8]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   134: begin
//row=9, col=6, rxregtablemod(row,col)=4243;
         wr_en_vec[8]=1;
         wr_address[8]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   135: begin
//row=9, col=7, rxregtablemod(row,col)=4275;
         wr_en_vec[8]=1;
         wr_address[8]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   136: begin
//row=9, col=8, rxregtablemod(row,col)=4307;
         wr_en_vec[8]=1;
         wr_address[8]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   137: begin
//row=9, col=9, rxregtablemod(row,col)=4339;
         wr_en_vec[8]=1;
         wr_address[8]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   138: begin
//row=9, col=10, rxregtablemod(row,col)=4371;
         wr_en_vec[8]=1;
         wr_address[8]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   139: begin
//row=9, col=11, rxregtablemod(row,col)=4403;
         wr_en_vec[8]=1;
         wr_address[8]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   140: begin
//row=9, col=12, rxregtablemod(row,col)=4435;
         wr_en_vec[8]=1;
         wr_address[8]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   141: begin
//row=9, col=13, rxregtablemod(row,col)=4467;
         wr_en_vec[8]=1;
         wr_address[8]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   142: begin
//row=9, col=14, rxregtablemod(row,col)=4499;
         wr_en_vec[8]=1;
         wr_address[8]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   143: begin
//row=9, col=15, rxregtablemod(row,col)=4531;
         wr_en_vec[8]=1;
         wr_address[8]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   144: begin
//row=9, col=16, rxregtablemod(row,col)=4563;
         wr_en_vec[8]=1;
         wr_address[8]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   145: begin
//row=10, col=1, rxregtablemod(row,col)=4595;
         wr_en_vec[9]=1;
         wr_address[9]=0;
//row=9, col=17, rxregtablemod(i,17)=4595;
         wr_en_vec[8]=1;
         wr_address[8]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   146: begin
//row=10, col=2, rxregtablemod(row,col)=4627;
         wr_en_vec[9]=1;
         wr_address[9]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   147: begin
//row=10, col=3, rxregtablemod(row,col)=4659;
         wr_en_vec[9]=1;
         wr_address[9]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   148: begin
//row=10, col=4, rxregtablemod(row,col)=4691;
         wr_en_vec[9]=1;
         wr_address[9]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   149: begin
//row=10, col=5, rxregtablemod(row,col)=4723;
         wr_en_vec[9]=1;
         wr_address[9]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   150: begin
//row=10, col=6, rxregtablemod(row,col)=4755;
         wr_en_vec[9]=1;
         wr_address[9]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   151: begin
//row=10, col=7, rxregtablemod(row,col)=4787;
         wr_en_vec[9]=1;
         wr_address[9]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   152: begin
//row=10, col=8, rxregtablemod(row,col)=4819;
         wr_en_vec[9]=1;
         wr_address[9]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   153: begin
//row=10, col=9, rxregtablemod(row,col)=4851;
         wr_en_vec[9]=1;
         wr_address[9]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   154: begin
//row=10, col=10, rxregtablemod(row,col)=4883;
         wr_en_vec[9]=1;
         wr_address[9]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   155: begin
//row=10, col=11, rxregtablemod(row,col)=4915;
         wr_en_vec[9]=1;
         wr_address[9]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   156: begin
//row=10, col=12, rxregtablemod(row,col)=4947;
         wr_en_vec[9]=1;
         wr_address[9]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   157: begin
//row=10, col=13, rxregtablemod(row,col)=4979;
         wr_en_vec[9]=1;
         wr_address[9]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   158: begin
//row=10, col=14, rxregtablemod(row,col)=5011;
         wr_en_vec[9]=1;
         wr_address[9]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   159: begin
//row=10, col=15, rxregtablemod(row,col)=5043;
         wr_en_vec[9]=1;
         wr_address[9]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   160: begin
//row=10, col=16, rxregtablemod(row,col)=5075;
         wr_en_vec[9]=1;
         wr_address[9]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   161: begin
//row=11, col=1, rxregtablemod(row,col)=5107;
         wr_en_vec[10]=1;
         wr_address[10]=0;
//row=10, col=17, rxregtablemod(i,17)=5107;
         wr_en_vec[9]=1;
         wr_address[9]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   162: begin
//row=11, col=2, rxregtablemod(row,col)=5139;
         wr_en_vec[10]=1;
         wr_address[10]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   163: begin
//row=11, col=3, rxregtablemod(row,col)=5171;
         wr_en_vec[10]=1;
         wr_address[10]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   164: begin
//row=11, col=4, rxregtablemod(row,col)=5203;
         wr_en_vec[10]=1;
         wr_address[10]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   165: begin
//row=11, col=5, rxregtablemod(row,col)=5235;
         wr_en_vec[10]=1;
         wr_address[10]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   166: begin
//row=11, col=6, rxregtablemod(row,col)=5267;
         wr_en_vec[10]=1;
         wr_address[10]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   167: begin
//row=11, col=7, rxregtablemod(row,col)=5299;
         wr_en_vec[10]=1;
         wr_address[10]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   168: begin
//row=11, col=8, rxregtablemod(row,col)=5331;
         wr_en_vec[10]=1;
         wr_address[10]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   169: begin
//row=11, col=9, rxregtablemod(row,col)=5363;
         wr_en_vec[10]=1;
         wr_address[10]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   170: begin
//row=11, col=10, rxregtablemod(row,col)=5395;
         wr_en_vec[10]=1;
         wr_address[10]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   171: begin
//row=11, col=11, rxregtablemod(row,col)=5427;
         wr_en_vec[10]=1;
         wr_address[10]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   172: begin
//row=11, col=12, rxregtablemod(row,col)=5459;
         wr_en_vec[10]=1;
         wr_address[10]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   173: begin
//row=11, col=13, rxregtablemod(row,col)=5491;
         wr_en_vec[10]=1;
         wr_address[10]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   174: begin
//row=11, col=14, rxregtablemod(row,col)=5523;
         wr_en_vec[10]=1;
         wr_address[10]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   175: begin
//row=11, col=15, rxregtablemod(row,col)=5555;
         wr_en_vec[10]=1;
         wr_address[10]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   176: begin
//row=11, col=16, rxregtablemod(row,col)=5587;
         wr_en_vec[10]=1;
         wr_address[10]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   177: begin
//row=12, col=1, rxregtablemod(row,col)=5619;
         wr_en_vec[11]=1;
         wr_address[11]=0;
//row=11, col=17, rxregtablemod(i,17)=5619;
         wr_en_vec[10]=1;
         wr_address[10]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   178: begin
//row=12, col=2, rxregtablemod(row,col)=5651;
         wr_en_vec[11]=1;
         wr_address[11]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   179: begin
//row=12, col=3, rxregtablemod(row,col)=5683;
         wr_en_vec[11]=1;
         wr_address[11]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   180: begin
//row=12, col=4, rxregtablemod(row,col)=5715;
         wr_en_vec[11]=1;
         wr_address[11]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   181: begin
//row=12, col=5, rxregtablemod(row,col)=5747;
         wr_en_vec[11]=1;
         wr_address[11]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   182: begin
//row=12, col=6, rxregtablemod(row,col)=5779;
         wr_en_vec[11]=1;
         wr_address[11]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   183: begin
//row=12, col=7, rxregtablemod(row,col)=5811;
         wr_en_vec[11]=1;
         wr_address[11]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   184: begin
//row=12, col=8, rxregtablemod(row,col)=5843;
         wr_en_vec[11]=1;
         wr_address[11]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   185: begin
//row=12, col=9, rxregtablemod(row,col)=5875;
         wr_en_vec[11]=1;
         wr_address[11]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   186: begin
//row=12, col=10, rxregtablemod(row,col)=5907;
         wr_en_vec[11]=1;
         wr_address[11]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   187: begin
//row=12, col=11, rxregtablemod(row,col)=5939;
         wr_en_vec[11]=1;
         wr_address[11]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   188: begin
//row=12, col=12, rxregtablemod(row,col)=5971;
         wr_en_vec[11]=1;
         wr_address[11]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   189: begin
//row=12, col=13, rxregtablemod(row,col)=6003;
         wr_en_vec[11]=1;
         wr_address[11]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   190: begin
//row=12, col=14, rxregtablemod(row,col)=6035;
         wr_en_vec[11]=1;
         wr_address[11]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   191: begin
//row=12, col=15, rxregtablemod(row,col)=6067;
         wr_en_vec[11]=1;
         wr_address[11]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   192: begin
//row=12, col=16, rxregtablemod(row,col)=6099;
         wr_en_vec[11]=1;
         wr_address[11]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   193: begin
//row=13, col=1, rxregtablemod(row,col)=6131;
         wr_en_vec[12]=1;
         wr_address[12]=0;
//row=12, col=17, rxregtablemod(i,17)=6131;
         wr_en_vec[11]=1;
         wr_address[11]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   194: begin
//row=13, col=2, rxregtablemod(row,col)=6163;
         wr_en_vec[12]=1;
         wr_address[12]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   195: begin
//row=13, col=3, rxregtablemod(row,col)=6195;
         wr_en_vec[12]=1;
         wr_address[12]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   196: begin
//row=13, col=4, rxregtablemod(row,col)=6227;
         wr_en_vec[12]=1;
         wr_address[12]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   197: begin
//row=13, col=5, rxregtablemod(row,col)=6259;
         wr_en_vec[12]=1;
         wr_address[12]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   198: begin
//row=13, col=6, rxregtablemod(row,col)=6291;
         wr_en_vec[12]=1;
         wr_address[12]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   199: begin
//row=13, col=7, rxregtablemod(row,col)=6323;
         wr_en_vec[12]=1;
         wr_address[12]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   200: begin
//row=13, col=8, rxregtablemod(row,col)=6355;
         wr_en_vec[12]=1;
         wr_address[12]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   201: begin
//row=13, col=9, rxregtablemod(row,col)=6387;
         wr_en_vec[12]=1;
         wr_address[12]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   202: begin
//row=13, col=10, rxregtablemod(row,col)=6419;
         wr_en_vec[12]=1;
         wr_address[12]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   203: begin
//row=13, col=11, rxregtablemod(row,col)=6451;
         wr_en_vec[12]=1;
         wr_address[12]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   204: begin
//row=13, col=12, rxregtablemod(row,col)=6483;
         wr_en_vec[12]=1;
         wr_address[12]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   205: begin
//row=13, col=13, rxregtablemod(row,col)=6515;
         wr_en_vec[12]=1;
         wr_address[12]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   206: begin
//row=13, col=14, rxregtablemod(row,col)=6547;
         wr_en_vec[12]=1;
         wr_address[12]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   207: begin
//row=13, col=15, rxregtablemod(row,col)=6579;
         wr_en_vec[12]=1;
         wr_address[12]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   208: begin
//row=13, col=16, rxregtablemod(row,col)=6611;
         wr_en_vec[12]=1;
         wr_address[12]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   209: begin
//row=14, col=1, rxregtablemod(row,col)=6643;
         wr_en_vec[13]=1;
         wr_address[13]=0;
//row=13, col=17, rxregtablemod(i,17)=6643;
         wr_en_vec[12]=1;
         wr_address[12]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   210: begin
//row=14, col=2, rxregtablemod(row,col)=6675;
         wr_en_vec[13]=1;
         wr_address[13]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   211: begin
//row=14, col=3, rxregtablemod(row,col)=6707;
         wr_en_vec[13]=1;
         wr_address[13]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   212: begin
//row=14, col=4, rxregtablemod(row,col)=6739;
         wr_en_vec[13]=1;
         wr_address[13]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   213: begin
//row=14, col=5, rxregtablemod(row,col)=6771;
         wr_en_vec[13]=1;
         wr_address[13]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   214: begin
//row=14, col=6, rxregtablemod(row,col)=6803;
         wr_en_vec[13]=1;
         wr_address[13]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   215: begin
//row=14, col=7, rxregtablemod(row,col)=6835;
         wr_en_vec[13]=1;
         wr_address[13]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   216: begin
//row=14, col=8, rxregtablemod(row,col)=6867;
         wr_en_vec[13]=1;
         wr_address[13]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   217: begin
//row=14, col=9, rxregtablemod(row,col)=6899;
         wr_en_vec[13]=1;
         wr_address[13]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   218: begin
//row=14, col=10, rxregtablemod(row,col)=6931;
         wr_en_vec[13]=1;
         wr_address[13]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   219: begin
//row=14, col=11, rxregtablemod(row,col)=6963;
         wr_en_vec[13]=1;
         wr_address[13]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   220: begin
//row=14, col=12, rxregtablemod(row,col)=6995;
         wr_en_vec[13]=1;
         wr_address[13]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   221: begin
//row=14, col=13, rxregtablemod(row,col)=7027;
         wr_en_vec[13]=1;
         wr_address[13]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   222: begin
//row=14, col=14, rxregtablemod(row,col)=7059;
         wr_en_vec[13]=1;
         wr_address[13]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   223: begin
//row=14, col=15, rxregtablemod(row,col)=7091;
         wr_en_vec[13]=1;
         wr_address[13]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   224: begin
//row=14, col=16, rxregtablemod(row,col)=7123;
         wr_en_vec[13]=1;
         wr_address[13]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   225: begin
//row=15, col=1, rxregtablemod(row,col)=7155;
         wr_en_vec[14]=1;
         wr_address[14]=0;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   226: begin
//row=15, col=2, rxregtablemod(row,col)=7187;
         wr_en_vec[14]=1;
         wr_address[14]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   227: begin
//row=15, col=3, rxregtablemod(row,col)=7219;
         wr_en_vec[14]=1;
         wr_address[14]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   228: begin
//row=15, col=4, rxregtablemod(row,col)=7251;
         wr_en_vec[14]=1;
         wr_address[14]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   229: begin
//row=15, col=5, rxregtablemod(row,col)=7283;
         wr_en_vec[14]=1;
         wr_address[14]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   230: begin
//row=15, col=6, rxregtablemod(row,col)=7315;
         wr_en_vec[14]=1;
         wr_address[14]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   231: begin
//row=15, col=7, rxregtablemod(row,col)=7347;
         wr_en_vec[14]=1;
         wr_address[14]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   232: begin
//row=15, col=8, rxregtablemod(row,col)=7379;
         wr_en_vec[14]=1;
         wr_address[14]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   233: begin
//row=15, col=9, rxregtablemod(row,col)=7411;
         wr_en_vec[14]=1;
         wr_address[14]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   234: begin
//row=15, col=10, rxregtablemod(row,col)=7443;
         wr_en_vec[14]=1;
         wr_address[14]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   235: begin
//row=15, col=11, rxregtablemod(row,col)=7475;
         wr_en_vec[14]=1;
         wr_address[14]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   236: begin
//row=15, col=12, rxregtablemod(row,col)=7507;
         wr_en_vec[14]=1;
         wr_address[14]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   237: begin
//row=15, col=13, rxregtablemod(row,col)=7539;
         wr_en_vec[14]=1;
         wr_address[14]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   238: begin
//row=15, col=14, rxregtablemod(row,col)=7571;
         wr_en_vec[14]=1;
         wr_address[14]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   239: begin
//row=15, col=15, rxregtablemod(row,col)=7603;
         wr_en_vec[14]=1;
         wr_address[14]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[15]=0;
         wr_address[15]=0;
       end
   240: begin
//row=16, col=1, rxregtablemod(row,col)=7635;
         wr_en_vec[15]=1;
         wr_address[15]=0;
//row=15, col=16, rxregtablemod(i,16)=7635;
         wr_en_vec[14]=1;
         wr_address[14]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
       end
   241: begin
//row=16, col=2, rxregtablemod(row,col)=7667;
         wr_en_vec[15]=1;
         wr_address[15]=1;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   242: begin
//row=16, col=3, rxregtablemod(row,col)=7699;
         wr_en_vec[15]=1;
         wr_address[15]=2;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   243: begin
//row=16, col=4, rxregtablemod(row,col)=7731;
         wr_en_vec[15]=1;
         wr_address[15]=3;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   244: begin
//row=16, col=5, rxregtablemod(row,col)=7763;
         wr_en_vec[15]=1;
         wr_address[15]=4;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   245: begin
//row=16, col=6, rxregtablemod(row,col)=7795;
         wr_en_vec[15]=1;
         wr_address[15]=5;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   246: begin
//row=16, col=7, rxregtablemod(row,col)=7827;
         wr_en_vec[15]=1;
         wr_address[15]=6;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   247: begin
//row=16, col=8, rxregtablemod(row,col)=7859;
         wr_en_vec[15]=1;
         wr_address[15]=7;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   248: begin
//row=16, col=9, rxregtablemod(row,col)=7891;
         wr_en_vec[15]=1;
         wr_address[15]=8;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   249: begin
//row=16, col=10, rxregtablemod(row,col)=7923;
         wr_en_vec[15]=1;
         wr_address[15]=9;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   250: begin
//row=16, col=11, rxregtablemod(row,col)=7955;
         wr_en_vec[15]=1;
         wr_address[15]=10;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   251: begin
//row=16, col=12, rxregtablemod(row,col)=7987;
         wr_en_vec[15]=1;
         wr_address[15]=11;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   252: begin
//row=16, col=13, rxregtablemod(row,col)=8019;
         wr_en_vec[15]=1;
         wr_address[15]=12;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   253: begin
//row=16, col=14, rxregtablemod(row,col)=8051;
         wr_en_vec[15]=1;
         wr_address[15]=13;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   254: begin
//row=16, col=15, rxregtablemod(row,col)=8083;
         wr_en_vec[15]=1;
         wr_address[15]=14;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   255: begin
//row=16, col=16, rxregtablemod(row,col)=8115;
         wr_en_vec[15]=1;
         wr_address[15]=15;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   256: begin
//row=16, col=17, rxregtablemod(row,col)=8147;
         wr_en_vec[15]=1;
         wr_address[15]=16;
         wr_en_vec[0]=0;
         wr_address[0]=0;
         wr_en_vec[1]=0;
         wr_address[1]=0;
         wr_en_vec[2]=0;
         wr_address[2]=0;
         wr_en_vec[3]=0;
         wr_address[3]=0;
         wr_en_vec[4]=0;
         wr_address[4]=0;
         wr_en_vec[5]=0;
         wr_address[5]=0;
         wr_en_vec[6]=0;
         wr_address[6]=0;
         wr_en_vec[7]=0;
         wr_address[7]=0;
         wr_en_vec[8]=0;
         wr_address[8]=0;
         wr_en_vec[9]=0;
         wr_address[9]=0;
         wr_en_vec[10]=0;
         wr_address[10]=0;
         wr_en_vec[11]=0;
         wr_address[11]=0;
         wr_en_vec[12]=0;
         wr_address[12]=0;
         wr_en_vec[13]=0;
         wr_address[13]=0;
         wr_en_vec[14]=0;
         wr_address[14]=0;
       end
   default: begin
              wr_en_vec[0]=0;
              wr_address[0]=0;
              wr_en_vec[1]=0;
              wr_address[1]=0;
              wr_en_vec[2]=0;
              wr_address[2]=0;
              wr_en_vec[3]=0;
              wr_address[3]=0;
              wr_en_vec[4]=0;
              wr_address[4]=0;
              wr_en_vec[5]=0;
              wr_address[5]=0;
              wr_en_vec[6]=0;
              wr_address[6]=0;
              wr_en_vec[7]=0;
              wr_address[7]=0;
              wr_en_vec[8]=0;
              wr_address[8]=0;
              wr_en_vec[9]=0;
              wr_address[9]=0;
              wr_en_vec[10]=0;
              wr_address[10]=0;
              wr_en_vec[11]=0;
              wr_address[11]=0;
              wr_en_vec[12]=0;
              wr_address[12]=0;
              wr_en_vec[13]=0;
              wr_address[13]=0;
              wr_en_vec[14]=0;
              wr_address[14]=0;
              wr_en_vec[15]=0;
              wr_address[15]=0;
            //first 64 ASM symbols of 0th cycle is skipped using this default case.
            end
  endcase
end
endmodule
