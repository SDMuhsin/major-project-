`timescale 1ns / 1ps

// Scripted from readselector_print.m 

module readselector_outputintf(outdata,rd_en_vec,rd_address_vec,memoutdata_vec,cyclecount,rd_en);
parameter ADDRESSWIDTH = 5;
parameter unloadMuxOutBits = 32;
parameter Kb = 14;//14*511=7154 systematic part

parameter CYCLECOUNTWIDTH = 8;//maxcycles=floor(7154/32)=223, width=ceil(log2(223))=8

output reg[unloadMuxOutBits-1:0] outdata;
output reg[Kb-1:0] rd_en_vec;
output [(Kb*ADDRESSWIDTH)-1:0] rd_address_vec;
input[(Kb*unloadMuxOutBits)-1:0] memoutdata_vec;
input[(CYCLECOUNTWIDTH)-1:0] cyclecount;
input rd_en;

reg[(ADDRESSWIDTH)-1:0] rd_address[Kb-1:0];
wire[(unloadMuxOutBits)-1:0] memoutdata[Kb-1:0];

genvar i;
generate
    for (i=0;i<Kb;i=i+1)begin:kb_loop
        assign rd_address_vec[ ((i+1)*ADDRESSWIDTH)-1:i*ADDRESSWIDTH]=rd_address[i];
        assign memoutdata[i]=memoutdata_vec[ ((i+1)*unloadMuxOutBits)-1:i*unloadMuxOutBits];
    end
endgenerate

always@(*) begin
  case(cyclecount)
   0: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   1: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=1;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   2: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=2;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   3: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=3;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   4: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=4;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   5: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=5;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   6: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=6;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   7: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=7;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   8: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=8;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   9: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=9;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   10: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=10;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   11: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=11;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   12: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=12;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   13: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=13;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   14: begin
         outdata=memoutdata[0];
         rd_en_vec[0]=rd_en;
         rd_address[0]=14;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   15: begin
         outdata={memoutdata[1][31:13],memoutdata[0][12:0]};
         rd_en_vec[0]=rd_en;
         rd_address[0]=15;
         rd_en_vec[1]=rd_en;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   16: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=1;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   17: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=2;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   18: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=3;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   19: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=4;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   20: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=5;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   21: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=6;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   22: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=7;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   23: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=8;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   24: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=9;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   25: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=10;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   26: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=11;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   27: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=12;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   28: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=13;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   29: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=14;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   30: begin
         outdata=memoutdata[1];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=15;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   31: begin
         outdata={memoutdata[2][31:12],memoutdata[1][11:0]};
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=rd_en;
         rd_address[1]=16;
         rd_en_vec[2]=rd_en;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   32: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=1;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   33: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=2;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   34: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=3;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   35: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=4;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   36: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=5;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   37: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=6;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   38: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=7;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   39: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=8;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   40: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=9;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   41: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=10;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   42: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=11;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   43: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=12;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   44: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=13;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   45: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=14;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   46: begin
         outdata=memoutdata[2];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=15;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   47: begin
         outdata={memoutdata[3][31:11],memoutdata[2][10:0]};
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=rd_en;
         rd_address[2]=16;
         rd_en_vec[3]=rd_en;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   48: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=1;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   49: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=2;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   50: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=3;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   51: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=4;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   52: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=5;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   53: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=6;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   54: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=7;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   55: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=8;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   56: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=9;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   57: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=10;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   58: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=11;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   59: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=12;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   60: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=13;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   61: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=14;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   62: begin
         outdata=memoutdata[3];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=15;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   63: begin
         outdata={memoutdata[4][31:10],memoutdata[3][9:0]};
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=rd_en;
         rd_address[3]=16;
         rd_en_vec[4]=rd_en;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   64: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=1;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   65: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=2;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   66: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=3;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   67: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=4;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   68: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=5;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   69: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=6;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   70: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=7;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   71: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=8;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   72: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=9;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   73: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=10;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   74: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=11;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   75: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=12;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   76: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=13;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   77: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=14;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   78: begin
         outdata=memoutdata[4];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=15;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   79: begin
         outdata={memoutdata[5][31:9],memoutdata[4][8:0]};
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=rd_en;
         rd_address[4]=16;
         rd_en_vec[5]=rd_en;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   80: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=1;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   81: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=2;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   82: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=3;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   83: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=4;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   84: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=5;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   85: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=6;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   86: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=7;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   87: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=8;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   88: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=9;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   89: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=10;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   90: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=11;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   91: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=12;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   92: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=13;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   93: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=14;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   94: begin
         outdata=memoutdata[5];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=15;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   95: begin
         outdata={memoutdata[6][31:8],memoutdata[5][7:0]};
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=rd_en;
         rd_address[5]=16;
         rd_en_vec[6]=rd_en;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   96: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=1;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   97: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=2;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   98: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=3;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   99: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=4;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   100: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=5;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   101: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=6;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   102: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=7;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   103: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=8;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   104: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=9;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   105: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=10;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   106: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=11;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   107: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=12;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   108: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=13;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   109: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=14;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   110: begin
         outdata=memoutdata[6];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=15;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   111: begin
         outdata={memoutdata[7][31:7],memoutdata[6][6:0]};
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=rd_en;
         rd_address[6]=16;
         rd_en_vec[7]=rd_en;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   112: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=1;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   113: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=2;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   114: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=3;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   115: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=4;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   116: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=5;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   117: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=6;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   118: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=7;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   119: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=8;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   120: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=9;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   121: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=10;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   122: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=11;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   123: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=12;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   124: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=13;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   125: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=14;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   126: begin
         outdata=memoutdata[7];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=15;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   127: begin
         outdata={memoutdata[8][31:6],memoutdata[7][5:0]};
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=rd_en;
         rd_address[7]=16;
         rd_en_vec[8]=rd_en;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   128: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=1;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   129: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=2;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   130: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=3;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   131: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=4;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   132: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=5;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   133: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=6;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   134: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=7;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   135: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=8;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   136: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=9;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   137: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=10;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   138: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=11;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   139: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=12;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   140: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=13;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   141: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=14;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   142: begin
         outdata=memoutdata[8];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=15;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   143: begin
         outdata={memoutdata[9][31:5],memoutdata[8][4:0]};
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=rd_en;
         rd_address[8]=16;
         rd_en_vec[9]=rd_en;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   144: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=1;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   145: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=2;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   146: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=3;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   147: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=4;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   148: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=5;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   149: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=6;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   150: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=7;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   151: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=8;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   152: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=9;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   153: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=10;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   154: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=11;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   155: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=12;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   156: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=13;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   157: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=14;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   158: begin
         outdata=memoutdata[9];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=15;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   159: begin
         outdata={memoutdata[10][31:4],memoutdata[9][3:0]};
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=rd_en;
         rd_address[9]=16;
         rd_en_vec[10]=rd_en;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   160: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=1;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   161: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=2;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   162: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=3;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   163: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=4;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   164: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=5;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   165: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=6;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   166: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=7;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   167: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=8;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   168: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=9;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   169: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=10;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   170: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=11;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   171: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=12;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   172: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=13;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   173: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=14;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   174: begin
         outdata=memoutdata[10];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=15;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   175: begin
         outdata={memoutdata[11][31:3],memoutdata[10][2:0]};
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=rd_en;
         rd_address[10]=16;
         rd_en_vec[11]=rd_en;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   176: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=1;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   177: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=2;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   178: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=3;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   179: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=4;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   180: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=5;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   181: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=6;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   182: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=7;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   183: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=8;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   184: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=9;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   185: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=10;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   186: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=11;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   187: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=12;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   188: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=13;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   189: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=14;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   190: begin
         outdata=memoutdata[11];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=15;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   191: begin
         outdata={memoutdata[12][31:2],memoutdata[11][1:0]};
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=rd_en;
         rd_address[11]=16;
         rd_en_vec[12]=rd_en;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   192: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=1;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   193: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=2;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   194: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=3;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   195: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=4;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   196: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=5;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   197: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=6;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   198: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=7;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   199: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=8;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   200: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=9;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   201: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=10;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   202: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=11;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   203: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=12;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   204: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=13;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   205: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=14;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   206: begin
         outdata=memoutdata[12];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=15;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
   207: begin
         outdata={memoutdata[13][31:1],memoutdata[12][0:0]};
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=rd_en;
         rd_address[12]=16;
         rd_en_vec[13]=rd_en;
         rd_address[13]=0;
       end
   208: begin
         outdata=memoutdata[13];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=1;
       end
   209: begin
         outdata=memoutdata[13];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=2;
       end
   210: begin
         outdata=memoutdata[13];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=3;
       end
   211: begin
         outdata=memoutdata[13];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=4;
       end
   212: begin
         outdata=memoutdata[13];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=5;
       end
   213: begin
         outdata=memoutdata[13];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=6;
       end
   214: begin
         outdata=memoutdata[13];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=7;
       end
   215: begin
         outdata=memoutdata[13];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=8;
       end
   216: begin
         outdata=memoutdata[13];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=9;
       end
   217: begin
         outdata=memoutdata[13];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=10;
       end
   218: begin
         outdata=memoutdata[13];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=11;
       end
   219: begin
         outdata=memoutdata[13];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=12;
       end
   220: begin
         outdata=memoutdata[13];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=13;
       end
   221: begin
         outdata=memoutdata[13];
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=14;
       end
   222: begin
         outdata={memoutdata[13][31:0]};
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=rd_en;
         rd_address[13]=15;
       end
   default: begin
         outdata=32'd0;
         rd_en_vec[0]=0;
         rd_address[0]=0;
         rd_en_vec[1]=0;
         rd_address[1]=0;
         rd_en_vec[2]=0;
         rd_address[2]=0;
         rd_en_vec[3]=0;
         rd_address[3]=0;
         rd_en_vec[4]=0;
         rd_address[4]=0;
         rd_en_vec[5]=0;
         rd_address[5]=0;
         rd_en_vec[6]=0;
         rd_address[6]=0;
         rd_en_vec[7]=0;
         rd_address[7]=0;
         rd_en_vec[8]=0;
         rd_address[8]=0;
         rd_en_vec[9]=0;
         rd_address[9]=0;
         rd_en_vec[10]=0;
         rd_address[10]=0;
         rd_en_vec[11]=0;
         rd_address[11]=0;
         rd_en_vec[12]=0;
         rd_address[12]=0;
         rd_en_vec[13]=0;
         rd_address[13]=0;
       end
  endcase
end//always
endmodule
