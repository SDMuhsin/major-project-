`timescale 1ns / 1ps
module LMem1To0_511_circ9_ys_yu_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        wr_en,
        feedback_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 15;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input [ADDRESSWIDTH-1:0]unloadAddress;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

input feedback_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        if(feedback_en) begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= fifoOut[i][c-1];
         end
        end
        else begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= ly0InConnector[i];
         end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
       0: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = fifoOut[1][11][w-1];
              unloadMuxOut[24] = fifoOut[2][11][w-1];
              unloadMuxOut[25] = fifoOut[3][11][w-1];
              unloadMuxOut[26] = fifoOut[4][11][w-1];
              unloadMuxOut[27] = fifoOut[5][11][w-1];
              unloadMuxOut[28] = fifoOut[6][11][w-1];
              unloadMuxOut[29] = fifoOut[7][11][w-1];
              unloadMuxOut[30] = fifoOut[8][11][w-1];
              unloadMuxOut[31] = fifoOut[9][11][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[10][11][w-1];
              unloadMuxOut[1] = fifoOut[11][11][w-1];
              unloadMuxOut[2] = fifoOut[12][11][w-1];
              unloadMuxOut[3] = fifoOut[13][11][w-1];
              unloadMuxOut[4] = fifoOut[14][11][w-1];
              unloadMuxOut[5] = fifoOut[15][11][w-1];
              unloadMuxOut[6] = fifoOut[16][11][w-1];
              unloadMuxOut[7] = fifoOut[17][11][w-1];
              unloadMuxOut[8] = fifoOut[18][11][w-1];
              unloadMuxOut[9] = fifoOut[19][11][w-1];
              unloadMuxOut[10] = fifoOut[20][11][w-1];
              unloadMuxOut[11] = fifoOut[21][11][w-1];
              unloadMuxOut[12] = fifoOut[22][11][w-1];
              unloadMuxOut[13] = fifoOut[23][11][w-1];
              unloadMuxOut[14] = fifoOut[24][11][w-1];
              unloadMuxOut[15] = fifoOut[25][11][w-1];
              unloadMuxOut[16] = fifoOut[0][10][w-1];
              unloadMuxOut[17] = fifoOut[1][10][w-1];
              unloadMuxOut[18] = fifoOut[2][10][w-1];
              unloadMuxOut[19] = fifoOut[3][10][w-1];
              unloadMuxOut[20] = fifoOut[4][10][w-1];
              unloadMuxOut[21] = fifoOut[5][10][w-1];
              unloadMuxOut[22] = fifoOut[6][10][w-1];
              unloadMuxOut[23] = fifoOut[7][10][w-1];
              unloadMuxOut[24] = fifoOut[8][10][w-1];
              unloadMuxOut[25] = fifoOut[9][10][w-1];
              unloadMuxOut[26] = fifoOut[10][10][w-1];
              unloadMuxOut[27] = fifoOut[11][10][w-1];
              unloadMuxOut[28] = fifoOut[12][10][w-1];
              unloadMuxOut[29] = fifoOut[13][10][w-1];
              unloadMuxOut[30] = fifoOut[14][10][w-1];
              unloadMuxOut[31] = fifoOut[15][10][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[16][10][w-1];
              unloadMuxOut[1] = fifoOut[17][10][w-1];
              unloadMuxOut[2] = fifoOut[18][10][w-1];
              unloadMuxOut[3] = fifoOut[19][10][w-1];
              unloadMuxOut[4] = fifoOut[20][10][w-1];
              unloadMuxOut[5] = fifoOut[21][10][w-1];
              unloadMuxOut[6] = fifoOut[22][10][w-1];
              unloadMuxOut[7] = fifoOut[23][10][w-1];
              unloadMuxOut[8] = fifoOut[24][10][w-1];
              unloadMuxOut[9] = fifoOut[25][10][w-1];
              unloadMuxOut[10] = fifoOut[0][9][w-1];
              unloadMuxOut[11] = fifoOut[1][9][w-1];
              unloadMuxOut[12] = fifoOut[2][9][w-1];
              unloadMuxOut[13] = fifoOut[3][9][w-1];
              unloadMuxOut[14] = fifoOut[4][9][w-1];
              unloadMuxOut[15] = fifoOut[5][9][w-1];
              unloadMuxOut[16] = fifoOut[6][9][w-1];
              unloadMuxOut[17] = fifoOut[7][9][w-1];
              unloadMuxOut[18] = fifoOut[8][9][w-1];
              unloadMuxOut[19] = fifoOut[9][9][w-1];
              unloadMuxOut[20] = fifoOut[10][9][w-1];
              unloadMuxOut[21] = fifoOut[11][9][w-1];
              unloadMuxOut[22] = fifoOut[12][9][w-1];
              unloadMuxOut[23] = fifoOut[13][9][w-1];
              unloadMuxOut[24] = fifoOut[14][9][w-1];
              unloadMuxOut[25] = fifoOut[15][9][w-1];
              unloadMuxOut[26] = fifoOut[16][9][w-1];
              unloadMuxOut[27] = fifoOut[17][9][w-1];
              unloadMuxOut[28] = fifoOut[18][9][w-1];
              unloadMuxOut[29] = fifoOut[26][14][w-1];
              unloadMuxOut[30] = fifoOut[27][14][w-1];
              unloadMuxOut[31] = fifoOut[28][14][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[29][14][w-1];
              unloadMuxOut[1] = fifoOut[30][14][w-1];
              unloadMuxOut[2] = fifoOut[31][14][w-1];
              unloadMuxOut[3] = fifoOut[32][14][w-1];
              unloadMuxOut[4] = fifoOut[33][14][w-1];
              unloadMuxOut[5] = fifoOut[34][14][w-1];
              unloadMuxOut[6] = fifoOut[35][14][w-1];
              unloadMuxOut[7] = fifoOut[36][14][w-1];
              unloadMuxOut[8] = fifoOut[37][14][w-1];
              unloadMuxOut[9] = fifoOut[38][14][w-1];
              unloadMuxOut[10] = fifoOut[39][14][w-1];
              unloadMuxOut[11] = fifoOut[40][14][w-1];
              unloadMuxOut[12] = fifoOut[41][14][w-1];
              unloadMuxOut[13] = fifoOut[42][14][w-1];
              unloadMuxOut[14] = fifoOut[43][14][w-1];
              unloadMuxOut[15] = fifoOut[44][14][w-1];
              unloadMuxOut[16] = fifoOut[45][14][w-1];
              unloadMuxOut[17] = fifoOut[46][14][w-1];
              unloadMuxOut[18] = fifoOut[47][14][w-1];
              unloadMuxOut[19] = fifoOut[48][14][w-1];
              unloadMuxOut[20] = fifoOut[49][14][w-1];
              unloadMuxOut[21] = fifoOut[50][14][w-1];
              unloadMuxOut[22] = fifoOut[51][14][w-1];
              unloadMuxOut[23] = fifoOut[26][13][w-1];
              unloadMuxOut[24] = fifoOut[27][13][w-1];
              unloadMuxOut[25] = fifoOut[28][13][w-1];
              unloadMuxOut[26] = fifoOut[29][13][w-1];
              unloadMuxOut[27] = fifoOut[30][13][w-1];
              unloadMuxOut[28] = fifoOut[31][13][w-1];
              unloadMuxOut[29] = fifoOut[32][13][w-1];
              unloadMuxOut[30] = fifoOut[33][13][w-1];
              unloadMuxOut[31] = fifoOut[34][13][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[35][13][w-1];
              unloadMuxOut[1] = fifoOut[36][13][w-1];
              unloadMuxOut[2] = fifoOut[37][13][w-1];
              unloadMuxOut[3] = fifoOut[38][13][w-1];
              unloadMuxOut[4] = fifoOut[39][13][w-1];
              unloadMuxOut[5] = fifoOut[40][13][w-1];
              unloadMuxOut[6] = fifoOut[41][13][w-1];
              unloadMuxOut[7] = fifoOut[42][13][w-1];
              unloadMuxOut[8] = fifoOut[43][13][w-1];
              unloadMuxOut[9] = fifoOut[44][13][w-1];
              unloadMuxOut[10] = fifoOut[45][13][w-1];
              unloadMuxOut[11] = fifoOut[46][13][w-1];
              unloadMuxOut[12] = fifoOut[47][13][w-1];
              unloadMuxOut[13] = fifoOut[48][13][w-1];
              unloadMuxOut[14] = fifoOut[49][13][w-1];
              unloadMuxOut[15] = fifoOut[50][13][w-1];
              unloadMuxOut[16] = fifoOut[51][13][w-1];
              unloadMuxOut[17] = fifoOut[26][12][w-1];
              unloadMuxOut[18] = fifoOut[27][12][w-1];
              unloadMuxOut[19] = fifoOut[28][12][w-1];
              unloadMuxOut[20] = fifoOut[29][12][w-1];
              unloadMuxOut[21] = fifoOut[30][12][w-1];
              unloadMuxOut[22] = fifoOut[31][12][w-1];
              unloadMuxOut[23] = fifoOut[32][12][w-1];
              unloadMuxOut[24] = fifoOut[33][12][w-1];
              unloadMuxOut[25] = fifoOut[34][12][w-1];
              unloadMuxOut[26] = fifoOut[35][12][w-1];
              unloadMuxOut[27] = fifoOut[36][12][w-1];
              unloadMuxOut[28] = fifoOut[37][12][w-1];
              unloadMuxOut[29] = fifoOut[38][12][w-1];
              unloadMuxOut[30] = fifoOut[39][12][w-1];
              unloadMuxOut[31] = fifoOut[40][12][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[41][12][w-1];
              unloadMuxOut[1] = fifoOut[42][12][w-1];
              unloadMuxOut[2] = fifoOut[43][12][w-1];
              unloadMuxOut[3] = fifoOut[44][12][w-1];
              unloadMuxOut[4] = fifoOut[45][12][w-1];
              unloadMuxOut[5] = fifoOut[46][12][w-1];
              unloadMuxOut[6] = fifoOut[47][12][w-1];
              unloadMuxOut[7] = fifoOut[48][12][w-1];
              unloadMuxOut[8] = fifoOut[49][12][w-1];
              unloadMuxOut[9] = fifoOut[50][12][w-1];
              unloadMuxOut[10] = fifoOut[51][12][w-1];
              unloadMuxOut[11] = fifoOut[26][11][w-1];
              unloadMuxOut[12] = fifoOut[27][11][w-1];
              unloadMuxOut[13] = fifoOut[28][11][w-1];
              unloadMuxOut[14] = fifoOut[29][11][w-1];
              unloadMuxOut[15] = fifoOut[30][11][w-1];
              unloadMuxOut[16] = fifoOut[31][11][w-1];
              unloadMuxOut[17] = fifoOut[32][11][w-1];
              unloadMuxOut[18] = fifoOut[33][11][w-1];
              unloadMuxOut[19] = fifoOut[34][11][w-1];
              unloadMuxOut[20] = fifoOut[35][11][w-1];
              unloadMuxOut[21] = fifoOut[36][11][w-1];
              unloadMuxOut[22] = fifoOut[37][11][w-1];
              unloadMuxOut[23] = fifoOut[38][11][w-1];
              unloadMuxOut[24] = fifoOut[39][11][w-1];
              unloadMuxOut[25] = fifoOut[40][11][w-1];
              unloadMuxOut[26] = fifoOut[41][11][w-1];
              unloadMuxOut[27] = fifoOut[42][11][w-1];
              unloadMuxOut[28] = fifoOut[43][11][w-1];
              unloadMuxOut[29] = fifoOut[44][11][w-1];
              unloadMuxOut[30] = fifoOut[45][11][w-1];
              unloadMuxOut[31] = fifoOut[46][11][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[47][11][w-1];
              unloadMuxOut[1] = fifoOut[48][11][w-1];
              unloadMuxOut[2] = fifoOut[49][11][w-1];
              unloadMuxOut[3] = fifoOut[50][11][w-1];
              unloadMuxOut[4] = fifoOut[51][11][w-1];
              unloadMuxOut[5] = fifoOut[26][10][w-1];
              unloadMuxOut[6] = fifoOut[27][10][w-1];
              unloadMuxOut[7] = fifoOut[28][10][w-1];
              unloadMuxOut[8] = fifoOut[29][10][w-1];
              unloadMuxOut[9] = fifoOut[30][10][w-1];
              unloadMuxOut[10] = fifoOut[31][10][w-1];
              unloadMuxOut[11] = fifoOut[32][10][w-1];
              unloadMuxOut[12] = fifoOut[33][10][w-1];
              unloadMuxOut[13] = fifoOut[34][10][w-1];
              unloadMuxOut[14] = fifoOut[35][10][w-1];
              unloadMuxOut[15] = fifoOut[36][10][w-1];
              unloadMuxOut[16] = fifoOut[37][10][w-1];
              unloadMuxOut[17] = fifoOut[38][10][w-1];
              unloadMuxOut[18] = fifoOut[39][10][w-1];
              unloadMuxOut[19] = fifoOut[40][10][w-1];
              unloadMuxOut[20] = fifoOut[41][10][w-1];
              unloadMuxOut[21] = fifoOut[42][10][w-1];
              unloadMuxOut[22] = fifoOut[43][10][w-1];
              unloadMuxOut[23] = fifoOut[44][10][w-1];
              unloadMuxOut[24] = fifoOut[45][10][w-1];
              unloadMuxOut[25] = fifoOut[46][10][w-1];
              unloadMuxOut[26] = fifoOut[47][10][w-1];
              unloadMuxOut[27] = fifoOut[48][10][w-1];
              unloadMuxOut[28] = fifoOut[49][10][w-1];
              unloadMuxOut[29] = fifoOut[50][10][w-1];
              unloadMuxOut[30] = fifoOut[51][10][w-1];
              unloadMuxOut[31] = fifoOut[26][9][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[27][9][w-1];
              unloadMuxOut[1] = fifoOut[28][9][w-1];
              unloadMuxOut[2] = fifoOut[29][9][w-1];
              unloadMuxOut[3] = fifoOut[30][9][w-1];
              unloadMuxOut[4] = fifoOut[31][9][w-1];
              unloadMuxOut[5] = fifoOut[32][9][w-1];
              unloadMuxOut[6] = fifoOut[33][9][w-1];
              unloadMuxOut[7] = fifoOut[34][9][w-1];
              unloadMuxOut[8] = fifoOut[35][9][w-1];
              unloadMuxOut[9] = fifoOut[36][9][w-1];
              unloadMuxOut[10] = fifoOut[37][9][w-1];
              unloadMuxOut[11] = fifoOut[38][9][w-1];
              unloadMuxOut[12] = fifoOut[39][9][w-1];
              unloadMuxOut[13] = fifoOut[40][9][w-1];
              unloadMuxOut[14] = fifoOut[41][9][w-1];
              unloadMuxOut[15] = fifoOut[42][9][w-1];
              unloadMuxOut[16] = fifoOut[43][9][w-1];
              unloadMuxOut[17] = fifoOut[44][9][w-1];
              unloadMuxOut[18] = fifoOut[45][9][w-1];
              unloadMuxOut[19] = fifoOut[46][9][w-1];
              unloadMuxOut[20] = fifoOut[47][9][w-1];
              unloadMuxOut[21] = fifoOut[48][9][w-1];
              unloadMuxOut[22] = fifoOut[49][9][w-1];
              unloadMuxOut[23] = fifoOut[50][9][w-1];
              unloadMuxOut[24] = fifoOut[51][9][w-1];
              unloadMuxOut[25] = fifoOut[26][8][w-1];
              unloadMuxOut[26] = fifoOut[27][8][w-1];
              unloadMuxOut[27] = fifoOut[28][8][w-1];
              unloadMuxOut[28] = fifoOut[29][8][w-1];
              unloadMuxOut[29] = fifoOut[30][8][w-1];
              unloadMuxOut[30] = fifoOut[31][8][w-1];
              unloadMuxOut[31] = fifoOut[32][8][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[33][8][w-1];
              unloadMuxOut[1] = fifoOut[34][8][w-1];
              unloadMuxOut[2] = fifoOut[35][8][w-1];
              unloadMuxOut[3] = fifoOut[36][8][w-1];
              unloadMuxOut[4] = fifoOut[37][8][w-1];
              unloadMuxOut[5] = fifoOut[38][8][w-1];
              unloadMuxOut[6] = fifoOut[39][8][w-1];
              unloadMuxOut[7] = fifoOut[40][8][w-1];
              unloadMuxOut[8] = fifoOut[41][8][w-1];
              unloadMuxOut[9] = fifoOut[42][8][w-1];
              unloadMuxOut[10] = fifoOut[43][8][w-1];
              unloadMuxOut[11] = fifoOut[44][8][w-1];
              unloadMuxOut[12] = fifoOut[45][8][w-1];
              unloadMuxOut[13] = fifoOut[46][8][w-1];
              unloadMuxOut[14] = fifoOut[47][8][w-1];
              unloadMuxOut[15] = fifoOut[48][8][w-1];
              unloadMuxOut[16] = fifoOut[49][8][w-1];
              unloadMuxOut[17] = fifoOut[50][8][w-1];
              unloadMuxOut[18] = fifoOut[51][8][w-1];
              unloadMuxOut[19] = fifoOut[26][7][w-1];
              unloadMuxOut[20] = fifoOut[27][7][w-1];
              unloadMuxOut[21] = fifoOut[28][7][w-1];
              unloadMuxOut[22] = fifoOut[29][7][w-1];
              unloadMuxOut[23] = fifoOut[30][7][w-1];
              unloadMuxOut[24] = fifoOut[31][7][w-1];
              unloadMuxOut[25] = fifoOut[32][7][w-1];
              unloadMuxOut[26] = fifoOut[33][7][w-1];
              unloadMuxOut[27] = fifoOut[34][7][w-1];
              unloadMuxOut[28] = fifoOut[35][7][w-1];
              unloadMuxOut[29] = fifoOut[36][7][w-1];
              unloadMuxOut[30] = fifoOut[37][7][w-1];
              unloadMuxOut[31] = fifoOut[38][7][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[39][7][w-1];
              unloadMuxOut[1] = fifoOut[40][7][w-1];
              unloadMuxOut[2] = fifoOut[41][7][w-1];
              unloadMuxOut[3] = fifoOut[42][7][w-1];
              unloadMuxOut[4] = fifoOut[43][7][w-1];
              unloadMuxOut[5] = fifoOut[44][7][w-1];
              unloadMuxOut[6] = fifoOut[45][7][w-1];
              unloadMuxOut[7] = fifoOut[46][7][w-1];
              unloadMuxOut[8] = fifoOut[47][7][w-1];
              unloadMuxOut[9] = fifoOut[48][7][w-1];
              unloadMuxOut[10] = fifoOut[49][7][w-1];
              unloadMuxOut[11] = fifoOut[50][7][w-1];
              unloadMuxOut[12] = fifoOut[51][7][w-1];
              unloadMuxOut[13] = fifoOut[26][6][w-1];
              unloadMuxOut[14] = fifoOut[27][6][w-1];
              unloadMuxOut[15] = fifoOut[28][6][w-1];
              unloadMuxOut[16] = fifoOut[29][6][w-1];
              unloadMuxOut[17] = fifoOut[30][6][w-1];
              unloadMuxOut[18] = fifoOut[31][6][w-1];
              unloadMuxOut[19] = fifoOut[32][6][w-1];
              unloadMuxOut[20] = fifoOut[33][6][w-1];
              unloadMuxOut[21] = fifoOut[34][6][w-1];
              unloadMuxOut[22] = fifoOut[35][6][w-1];
              unloadMuxOut[23] = fifoOut[36][6][w-1];
              unloadMuxOut[24] = fifoOut[37][6][w-1];
              unloadMuxOut[25] = fifoOut[38][6][w-1];
              unloadMuxOut[26] = fifoOut[39][6][w-1];
              unloadMuxOut[27] = fifoOut[40][6][w-1];
              unloadMuxOut[28] = fifoOut[41][6][w-1];
              unloadMuxOut[29] = fifoOut[42][6][w-1];
              unloadMuxOut[30] = fifoOut[43][6][w-1];
              unloadMuxOut[31] = fifoOut[44][6][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[45][6][w-1];
              unloadMuxOut[1] = fifoOut[46][6][w-1];
              unloadMuxOut[2] = fifoOut[47][6][w-1];
              unloadMuxOut[3] = fifoOut[48][6][w-1];
              unloadMuxOut[4] = fifoOut[49][6][w-1];
              unloadMuxOut[5] = fifoOut[50][6][w-1];
              unloadMuxOut[6] = fifoOut[51][6][w-1];
              unloadMuxOut[7] = fifoOut[26][5][w-1];
              unloadMuxOut[8] = fifoOut[27][5][w-1];
              unloadMuxOut[9] = fifoOut[28][5][w-1];
              unloadMuxOut[10] = fifoOut[29][5][w-1];
              unloadMuxOut[11] = fifoOut[30][5][w-1];
              unloadMuxOut[12] = fifoOut[31][5][w-1];
              unloadMuxOut[13] = fifoOut[32][5][w-1];
              unloadMuxOut[14] = fifoOut[33][5][w-1];
              unloadMuxOut[15] = fifoOut[34][5][w-1];
              unloadMuxOut[16] = fifoOut[35][5][w-1];
              unloadMuxOut[17] = fifoOut[36][5][w-1];
              unloadMuxOut[18] = fifoOut[37][5][w-1];
              unloadMuxOut[19] = fifoOut[38][5][w-1];
              unloadMuxOut[20] = fifoOut[39][5][w-1];
              unloadMuxOut[21] = fifoOut[40][5][w-1];
              unloadMuxOut[22] = fifoOut[41][5][w-1];
              unloadMuxOut[23] = fifoOut[42][5][w-1];
              unloadMuxOut[24] = fifoOut[43][5][w-1];
              unloadMuxOut[25] = fifoOut[44][5][w-1];
              unloadMuxOut[26] = fifoOut[45][5][w-1];
              unloadMuxOut[27] = fifoOut[46][5][w-1];
              unloadMuxOut[28] = fifoOut[47][5][w-1];
              unloadMuxOut[29] = fifoOut[48][5][w-1];
              unloadMuxOut[30] = fifoOut[49][5][w-1];
              unloadMuxOut[31] = fifoOut[50][5][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[51][5][w-1];
              unloadMuxOut[1] = fifoOut[26][4][w-1];
              unloadMuxOut[2] = fifoOut[27][4][w-1];
              unloadMuxOut[3] = fifoOut[28][4][w-1];
              unloadMuxOut[4] = fifoOut[29][4][w-1];
              unloadMuxOut[5] = fifoOut[30][4][w-1];
              unloadMuxOut[6] = fifoOut[31][4][w-1];
              unloadMuxOut[7] = fifoOut[32][4][w-1];
              unloadMuxOut[8] = fifoOut[33][4][w-1];
              unloadMuxOut[9] = fifoOut[34][4][w-1];
              unloadMuxOut[10] = fifoOut[35][4][w-1];
              unloadMuxOut[11] = fifoOut[36][4][w-1];
              unloadMuxOut[12] = fifoOut[37][4][w-1];
              unloadMuxOut[13] = fifoOut[38][4][w-1];
              unloadMuxOut[14] = fifoOut[39][4][w-1];
              unloadMuxOut[15] = fifoOut[40][4][w-1];
              unloadMuxOut[16] = fifoOut[41][4][w-1];
              unloadMuxOut[17] = fifoOut[42][4][w-1];
              unloadMuxOut[18] = fifoOut[43][4][w-1];
              unloadMuxOut[19] = fifoOut[44][4][w-1];
              unloadMuxOut[20] = fifoOut[45][4][w-1];
              unloadMuxOut[21] = fifoOut[46][4][w-1];
              unloadMuxOut[22] = fifoOut[47][4][w-1];
              unloadMuxOut[23] = fifoOut[48][4][w-1];
              unloadMuxOut[24] = fifoOut[49][4][w-1];
              unloadMuxOut[25] = fifoOut[50][4][w-1];
              unloadMuxOut[26] = fifoOut[51][4][w-1];
              unloadMuxOut[27] = fifoOut[26][3][w-1];
              unloadMuxOut[28] = fifoOut[27][3][w-1];
              unloadMuxOut[29] = fifoOut[28][3][w-1];
              unloadMuxOut[30] = fifoOut[29][3][w-1];
              unloadMuxOut[31] = fifoOut[30][3][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[31][3][w-1];
              unloadMuxOut[1] = fifoOut[32][3][w-1];
              unloadMuxOut[2] = fifoOut[33][3][w-1];
              unloadMuxOut[3] = fifoOut[34][3][w-1];
              unloadMuxOut[4] = fifoOut[35][3][w-1];
              unloadMuxOut[5] = fifoOut[36][3][w-1];
              unloadMuxOut[6] = fifoOut[37][3][w-1];
              unloadMuxOut[7] = fifoOut[38][3][w-1];
              unloadMuxOut[8] = fifoOut[39][3][w-1];
              unloadMuxOut[9] = fifoOut[40][3][w-1];
              unloadMuxOut[10] = fifoOut[41][3][w-1];
              unloadMuxOut[11] = fifoOut[42][3][w-1];
              unloadMuxOut[12] = fifoOut[43][3][w-1];
              unloadMuxOut[13] = fifoOut[44][3][w-1];
              unloadMuxOut[14] = fifoOut[45][3][w-1];
              unloadMuxOut[15] = fifoOut[46][3][w-1];
              unloadMuxOut[16] = fifoOut[47][3][w-1];
              unloadMuxOut[17] = fifoOut[48][3][w-1];
              unloadMuxOut[18] = fifoOut[49][3][w-1];
              unloadMuxOut[19] = fifoOut[50][3][w-1];
              unloadMuxOut[20] = fifoOut[51][3][w-1];
              unloadMuxOut[21] = fifoOut[26][2][w-1];
              unloadMuxOut[22] = fifoOut[27][2][w-1];
              unloadMuxOut[23] = fifoOut[28][2][w-1];
              unloadMuxOut[24] = fifoOut[29][2][w-1];
              unloadMuxOut[25] = fifoOut[30][2][w-1];
              unloadMuxOut[26] = fifoOut[31][2][w-1];
              unloadMuxOut[27] = fifoOut[32][2][w-1];
              unloadMuxOut[28] = fifoOut[33][2][w-1];
              unloadMuxOut[29] = fifoOut[34][2][w-1];
              unloadMuxOut[30] = fifoOut[35][2][w-1];
              unloadMuxOut[31] = fifoOut[36][2][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[37][2][w-1];
              unloadMuxOut[1] = fifoOut[38][2][w-1];
              unloadMuxOut[2] = fifoOut[39][2][w-1];
              unloadMuxOut[3] = fifoOut[40][2][w-1];
              unloadMuxOut[4] = fifoOut[41][2][w-1];
              unloadMuxOut[5] = fifoOut[42][2][w-1];
              unloadMuxOut[6] = fifoOut[43][2][w-1];
              unloadMuxOut[7] = fifoOut[44][2][w-1];
              unloadMuxOut[8] = fifoOut[45][2][w-1];
              unloadMuxOut[9] = fifoOut[46][2][w-1];
              unloadMuxOut[10] = fifoOut[47][2][w-1];
              unloadMuxOut[11] = fifoOut[48][2][w-1];
              unloadMuxOut[12] = fifoOut[49][2][w-1];
              unloadMuxOut[13] = fifoOut[50][2][w-1];
              unloadMuxOut[14] = fifoOut[51][2][w-1];
              unloadMuxOut[15] = fifoOut[26][1][w-1];
              unloadMuxOut[16] = fifoOut[27][1][w-1];
              unloadMuxOut[17] = fifoOut[28][1][w-1];
              unloadMuxOut[18] = fifoOut[29][1][w-1];
              unloadMuxOut[19] = fifoOut[30][1][w-1];
              unloadMuxOut[20] = fifoOut[31][1][w-1];
              unloadMuxOut[21] = fifoOut[32][1][w-1];
              unloadMuxOut[22] = fifoOut[33][1][w-1];
              unloadMuxOut[23] = fifoOut[34][1][w-1];
              unloadMuxOut[24] = fifoOut[35][1][w-1];
              unloadMuxOut[25] = fifoOut[36][1][w-1];
              unloadMuxOut[26] = fifoOut[37][1][w-1];
              unloadMuxOut[27] = fifoOut[38][1][w-1];
              unloadMuxOut[28] = fifoOut[39][1][w-1];
              unloadMuxOut[29] = fifoOut[40][1][w-1];
              unloadMuxOut[30] = fifoOut[41][1][w-1];
              unloadMuxOut[31] = fifoOut[42][1][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[43][1][w-1];
              unloadMuxOut[1] = fifoOut[44][1][w-1];
              unloadMuxOut[2] = fifoOut[45][1][w-1];
              unloadMuxOut[3] = fifoOut[46][1][w-1];
              unloadMuxOut[4] = fifoOut[47][1][w-1];
              unloadMuxOut[5] = fifoOut[48][1][w-1];
              unloadMuxOut[6] = fifoOut[49][1][w-1];
              unloadMuxOut[7] = fifoOut[0][14][w-1];
              unloadMuxOut[8] = fifoOut[1][14][w-1];
              unloadMuxOut[9] = fifoOut[2][14][w-1];
              unloadMuxOut[10] = fifoOut[3][14][w-1];
              unloadMuxOut[11] = fifoOut[4][14][w-1];
              unloadMuxOut[12] = fifoOut[5][14][w-1];
              unloadMuxOut[13] = fifoOut[6][14][w-1];
              unloadMuxOut[14] = fifoOut[7][14][w-1];
              unloadMuxOut[15] = fifoOut[8][14][w-1];
              unloadMuxOut[16] = fifoOut[9][14][w-1];
              unloadMuxOut[17] = fifoOut[10][14][w-1];
              unloadMuxOut[18] = fifoOut[11][14][w-1];
              unloadMuxOut[19] = fifoOut[12][14][w-1];
              unloadMuxOut[20] = fifoOut[13][14][w-1];
              unloadMuxOut[21] = fifoOut[14][14][w-1];
              unloadMuxOut[22] = fifoOut[15][14][w-1];
              unloadMuxOut[23] = fifoOut[16][14][w-1];
              unloadMuxOut[24] = fifoOut[17][14][w-1];
              unloadMuxOut[25] = fifoOut[18][14][w-1];
              unloadMuxOut[26] = fifoOut[19][14][w-1];
              unloadMuxOut[27] = fifoOut[20][14][w-1];
              unloadMuxOut[28] = fifoOut[21][14][w-1];
              unloadMuxOut[29] = fifoOut[22][14][w-1];
              unloadMuxOut[30] = fifoOut[23][14][w-1];
              unloadMuxOut[31] = fifoOut[24][14][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[25][14][w-1];
              unloadMuxOut[1] = fifoOut[0][13][w-1];
              unloadMuxOut[2] = fifoOut[1][13][w-1];
              unloadMuxOut[3] = fifoOut[2][13][w-1];
              unloadMuxOut[4] = fifoOut[3][13][w-1];
              unloadMuxOut[5] = fifoOut[4][13][w-1];
              unloadMuxOut[6] = fifoOut[5][13][w-1];
              unloadMuxOut[7] = fifoOut[6][13][w-1];
              unloadMuxOut[8] = fifoOut[7][13][w-1];
              unloadMuxOut[9] = fifoOut[8][13][w-1];
              unloadMuxOut[10] = fifoOut[9][13][w-1];
              unloadMuxOut[11] = fifoOut[10][13][w-1];
              unloadMuxOut[12] = fifoOut[11][13][w-1];
              unloadMuxOut[13] = fifoOut[12][13][w-1];
              unloadMuxOut[14] = fifoOut[13][13][w-1];
              unloadMuxOut[15] = fifoOut[14][13][w-1];
              unloadMuxOut[16] = fifoOut[15][13][w-1];
              unloadMuxOut[17] = fifoOut[16][13][w-1];
              unloadMuxOut[18] = fifoOut[17][13][w-1];
              unloadMuxOut[19] = fifoOut[18][13][w-1];
              unloadMuxOut[20] = fifoOut[19][13][w-1];
              unloadMuxOut[21] = fifoOut[20][13][w-1];
              unloadMuxOut[22] = fifoOut[21][13][w-1];
              unloadMuxOut[23] = fifoOut[22][13][w-1];
              unloadMuxOut[24] = fifoOut[23][13][w-1];
              unloadMuxOut[25] = fifoOut[24][13][w-1];
              unloadMuxOut[26] = fifoOut[25][13][w-1];
              unloadMuxOut[27] = fifoOut[0][12][w-1];
              unloadMuxOut[28] = fifoOut[1][12][w-1];
              unloadMuxOut[29] = fifoOut[2][12][w-1];
              unloadMuxOut[30] = fifoOut[3][12][w-1];
              unloadMuxOut[31] = fifoOut[4][12][w-1];
       end
       16: begin
              unloadMuxOut[0] = fifoOut[5][12][w-1];
              unloadMuxOut[1] = fifoOut[6][12][w-1];
              unloadMuxOut[2] = fifoOut[7][12][w-1];
              unloadMuxOut[3] = fifoOut[8][12][w-1];
              unloadMuxOut[4] = fifoOut[9][12][w-1];
              unloadMuxOut[5] = fifoOut[10][12][w-1];
              unloadMuxOut[6] = fifoOut[11][12][w-1];
              unloadMuxOut[7] = fifoOut[12][12][w-1];
              unloadMuxOut[8] = fifoOut[13][12][w-1];
              unloadMuxOut[9] = fifoOut[14][12][w-1];
              unloadMuxOut[10] = fifoOut[15][12][w-1];
              unloadMuxOut[11] = fifoOut[16][12][w-1];
              unloadMuxOut[12] = fifoOut[17][12][w-1];
              unloadMuxOut[13] = fifoOut[18][12][w-1];
              unloadMuxOut[14] = fifoOut[19][12][w-1];
              unloadMuxOut[15] = fifoOut[20][12][w-1];
              unloadMuxOut[16] = fifoOut[21][12][w-1];
              unloadMuxOut[17] = fifoOut[22][12][w-1];
              unloadMuxOut[18] = fifoOut[23][12][w-1];
              unloadMuxOut[19] = fifoOut[24][12][w-1];
              unloadMuxOut[20] = fifoOut[25][12][w-1];
              unloadMuxOut[21] = fifoOut[0][11][w-1];
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0;
             end
       end
    endcase
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[43][4];
              muxOutConnector[45] = fifoOut[44][4];
              muxOutConnector[46] = fifoOut[45][4];
              muxOutConnector[47] = fifoOut[46][4];
              muxOutConnector[48] = fifoOut[47][4];
              muxOutConnector[49] = fifoOut[48][4];
              muxOutConnector[50] = fifoOut[49][4];
              muxOutConnector[51] = fifoOut[50][4];
       end
       1: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[43][4];
              muxOutConnector[45] = fifoOut[44][4];
              muxOutConnector[46] = fifoOut[45][4];
              muxOutConnector[47] = fifoOut[46][4];
              muxOutConnector[48] = fifoOut[47][4];
              muxOutConnector[49] = fifoOut[48][4];
              muxOutConnector[50] = fifoOut[49][4];
              muxOutConnector[51] = fifoOut[50][4];
       end
       2: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[43][4];
              muxOutConnector[45] = fifoOut[44][4];
              muxOutConnector[46] = fifoOut[45][4];
              muxOutConnector[47] = fifoOut[46][4];
              muxOutConnector[48] = fifoOut[47][4];
              muxOutConnector[49] = fifoOut[48][4];
              muxOutConnector[50] = fifoOut[49][4];
              muxOutConnector[51] = fifoOut[50][4];
       end
       3: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[43][4];
              muxOutConnector[45] = fifoOut[44][4];
              muxOutConnector[46] = fifoOut[45][4];
              muxOutConnector[47] = fifoOut[46][4];
              muxOutConnector[48] = fifoOut[47][4];
              muxOutConnector[49] = fifoOut[48][4];
              muxOutConnector[50] = fifoOut[49][4];
              muxOutConnector[51] = fifoOut[50][4];
       end
       4: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[19][3];
              muxOutConnector[45] = fifoOut[20][3];
              muxOutConnector[46] = fifoOut[21][3];
              muxOutConnector[47] = fifoOut[22][3];
              muxOutConnector[48] = fifoOut[23][3];
              muxOutConnector[49] = fifoOut[24][3];
              muxOutConnector[50] = fifoOut[25][3];
              muxOutConnector[51] = fifoOut[0][2];
       end
       5: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][3];
              muxOutConnector[27] = fifoOut[2][3];
              muxOutConnector[28] = fifoOut[3][3];
              muxOutConnector[29] = fifoOut[4][3];
              muxOutConnector[30] = fifoOut[5][3];
              muxOutConnector[31] = fifoOut[6][3];
              muxOutConnector[32] = fifoOut[7][3];
              muxOutConnector[33] = fifoOut[8][3];
              muxOutConnector[34] = fifoOut[9][3];
              muxOutConnector[35] = fifoOut[10][3];
              muxOutConnector[36] = fifoOut[11][3];
              muxOutConnector[37] = fifoOut[12][3];
              muxOutConnector[38] = fifoOut[13][3];
              muxOutConnector[39] = fifoOut[14][3];
              muxOutConnector[40] = fifoOut[15][3];
              muxOutConnector[41] = fifoOut[16][3];
              muxOutConnector[42] = fifoOut[17][3];
              muxOutConnector[43] = fifoOut[18][3];
              muxOutConnector[44] = fifoOut[19][3];
              muxOutConnector[45] = fifoOut[20][3];
              muxOutConnector[46] = fifoOut[21][3];
              muxOutConnector[47] = fifoOut[22][3];
              muxOutConnector[48] = fifoOut[23][3];
              muxOutConnector[49] = fifoOut[24][3];
              muxOutConnector[50] = fifoOut[25][3];
              muxOutConnector[51] = fifoOut[0][2];
       end
       6: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][3];
              muxOutConnector[27] = fifoOut[2][3];
              muxOutConnector[28] = fifoOut[3][3];
              muxOutConnector[29] = fifoOut[4][3];
              muxOutConnector[30] = fifoOut[5][3];
              muxOutConnector[31] = fifoOut[6][3];
              muxOutConnector[32] = fifoOut[7][3];
              muxOutConnector[33] = fifoOut[8][3];
              muxOutConnector[34] = fifoOut[9][3];
              muxOutConnector[35] = fifoOut[10][3];
              muxOutConnector[36] = fifoOut[11][3];
              muxOutConnector[37] = fifoOut[12][3];
              muxOutConnector[38] = fifoOut[13][3];
              muxOutConnector[39] = fifoOut[14][3];
              muxOutConnector[40] = fifoOut[15][3];
              muxOutConnector[41] = fifoOut[16][3];
              muxOutConnector[42] = fifoOut[17][3];
              muxOutConnector[43] = fifoOut[18][3];
              muxOutConnector[44] = fifoOut[19][3];
              muxOutConnector[45] = fifoOut[20][3];
              muxOutConnector[46] = fifoOut[21][3];
              muxOutConnector[47] = fifoOut[22][3];
              muxOutConnector[48] = fifoOut[23][3];
              muxOutConnector[49] = fifoOut[24][3];
              muxOutConnector[50] = fifoOut[25][3];
              muxOutConnector[51] = fifoOut[0][2];
       end
       7: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][3];
              muxOutConnector[27] = fifoOut[2][3];
              muxOutConnector[28] = fifoOut[3][3];
              muxOutConnector[29] = fifoOut[4][3];
              muxOutConnector[30] = fifoOut[5][3];
              muxOutConnector[31] = fifoOut[6][3];
              muxOutConnector[32] = fifoOut[7][3];
              muxOutConnector[33] = fifoOut[8][3];
              muxOutConnector[34] = fifoOut[9][3];
              muxOutConnector[35] = fifoOut[10][3];
              muxOutConnector[36] = fifoOut[11][3];
              muxOutConnector[37] = fifoOut[12][3];
              muxOutConnector[38] = fifoOut[13][3];
              muxOutConnector[39] = fifoOut[14][3];
              muxOutConnector[40] = fifoOut[15][3];
              muxOutConnector[41] = fifoOut[16][3];
              muxOutConnector[42] = fifoOut[17][3];
              muxOutConnector[43] = fifoOut[18][3];
              muxOutConnector[44] = fifoOut[19][3];
              muxOutConnector[45] = fifoOut[20][3];
              muxOutConnector[46] = fifoOut[21][3];
              muxOutConnector[47] = fifoOut[22][3];
              muxOutConnector[48] = fifoOut[23][3];
              muxOutConnector[49] = fifoOut[24][3];
              muxOutConnector[50] = fifoOut[25][3];
              muxOutConnector[51] = fifoOut[0][2];
       end
       8: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][3];
              muxOutConnector[27] = fifoOut[2][3];
              muxOutConnector[28] = fifoOut[3][3];
              muxOutConnector[29] = fifoOut[4][3];
              muxOutConnector[30] = fifoOut[5][3];
              muxOutConnector[31] = fifoOut[6][3];
              muxOutConnector[32] = fifoOut[7][3];
              muxOutConnector[33] = fifoOut[8][3];
              muxOutConnector[34] = fifoOut[9][3];
              muxOutConnector[35] = fifoOut[10][3];
              muxOutConnector[36] = fifoOut[11][3];
              muxOutConnector[37] = fifoOut[12][3];
              muxOutConnector[38] = fifoOut[13][3];
              muxOutConnector[39] = fifoOut[14][3];
              muxOutConnector[40] = fifoOut[15][3];
              muxOutConnector[41] = fifoOut[16][3];
              muxOutConnector[42] = fifoOut[17][3];
              muxOutConnector[43] = fifoOut[18][3];
              muxOutConnector[44] = fifoOut[19][3];
              muxOutConnector[45] = fifoOut[20][3];
              muxOutConnector[46] = fifoOut[21][3];
              muxOutConnector[47] = fifoOut[22][3];
              muxOutConnector[48] = fifoOut[23][3];
              muxOutConnector[49] = fifoOut[24][3];
              muxOutConnector[50] = fifoOut[25][3];
              muxOutConnector[51] = fifoOut[0][2];
       end
       9: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[50][0];
              muxOutConnector[16] = fifoOut[51][0];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][3];
              muxOutConnector[27] = fifoOut[2][3];
              muxOutConnector[28] = fifoOut[3][3];
              muxOutConnector[29] = fifoOut[4][3];
              muxOutConnector[30] = fifoOut[5][3];
              muxOutConnector[31] = fifoOut[6][3];
              muxOutConnector[32] = fifoOut[7][3];
              muxOutConnector[33] = fifoOut[8][3];
              muxOutConnector[34] = fifoOut[9][3];
              muxOutConnector[35] = fifoOut[10][3];
              muxOutConnector[36] = fifoOut[11][3];
              muxOutConnector[37] = fifoOut[12][3];
              muxOutConnector[38] = fifoOut[13][3];
              muxOutConnector[39] = fifoOut[14][3];
              muxOutConnector[40] = fifoOut[15][3];
              muxOutConnector[41] = fifoOut[16][3];
              muxOutConnector[42] = fifoOut[17][3];
              muxOutConnector[43] = fifoOut[18][3];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       10: begin
              muxOutConnector[0] = fifoOut[35][0];
              muxOutConnector[1] = fifoOut[36][0];
              muxOutConnector[2] = fifoOut[37][0];
              muxOutConnector[3] = fifoOut[38][0];
              muxOutConnector[4] = fifoOut[39][0];
              muxOutConnector[5] = fifoOut[40][0];
              muxOutConnector[6] = fifoOut[41][0];
              muxOutConnector[7] = fifoOut[42][0];
              muxOutConnector[8] = fifoOut[43][0];
              muxOutConnector[9] = fifoOut[44][0];
              muxOutConnector[10] = fifoOut[45][0];
              muxOutConnector[11] = fifoOut[46][0];
              muxOutConnector[12] = fifoOut[47][0];
              muxOutConnector[13] = fifoOut[48][0];
              muxOutConnector[14] = fifoOut[49][0];
              muxOutConnector[15] = fifoOut[50][0];
              muxOutConnector[16] = fifoOut[51][0];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       11: begin
              muxOutConnector[0] = fifoOut[35][0];
              muxOutConnector[1] = fifoOut[36][0];
              muxOutConnector[2] = fifoOut[37][0];
              muxOutConnector[3] = fifoOut[38][0];
              muxOutConnector[4] = fifoOut[39][0];
              muxOutConnector[5] = fifoOut[40][0];
              muxOutConnector[6] = fifoOut[41][0];
              muxOutConnector[7] = fifoOut[42][0];
              muxOutConnector[8] = fifoOut[43][0];
              muxOutConnector[9] = fifoOut[44][0];
              muxOutConnector[10] = fifoOut[45][0];
              muxOutConnector[11] = fifoOut[46][0];
              muxOutConnector[12] = fifoOut[47][0];
              muxOutConnector[13] = fifoOut[48][0];
              muxOutConnector[14] = fifoOut[49][0];
              muxOutConnector[15] = fifoOut[50][0];
              muxOutConnector[16] = fifoOut[51][0];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       12: begin
              muxOutConnector[0] = fifoOut[35][0];
              muxOutConnector[1] = fifoOut[36][0];
              muxOutConnector[2] = fifoOut[37][0];
              muxOutConnector[3] = fifoOut[38][0];
              muxOutConnector[4] = fifoOut[39][0];
              muxOutConnector[5] = fifoOut[40][0];
              muxOutConnector[6] = fifoOut[41][0];
              muxOutConnector[7] = fifoOut[42][0];
              muxOutConnector[8] = fifoOut[43][0];
              muxOutConnector[9] = fifoOut[44][0];
              muxOutConnector[10] = fifoOut[45][0];
              muxOutConnector[11] = fifoOut[46][0];
              muxOutConnector[12] = fifoOut[47][0];
              muxOutConnector[13] = fifoOut[48][0];
              muxOutConnector[14] = fifoOut[49][0];
              muxOutConnector[15] = fifoOut[50][0];
              muxOutConnector[16] = fifoOut[51][0];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       13: begin
              muxOutConnector[0] = fifoOut[35][0];
              muxOutConnector[1] = fifoOut[36][0];
              muxOutConnector[2] = fifoOut[37][0];
              muxOutConnector[3] = fifoOut[38][0];
              muxOutConnector[4] = fifoOut[39][0];
              muxOutConnector[5] = fifoOut[40][0];
              muxOutConnector[6] = fifoOut[41][0];
              muxOutConnector[7] = fifoOut[42][0];
              muxOutConnector[8] = fifoOut[43][0];
              muxOutConnector[9] = fifoOut[44][0];
              muxOutConnector[10] = fifoOut[45][0];
              muxOutConnector[11] = fifoOut[46][0];
              muxOutConnector[12] = fifoOut[47][0];
              muxOutConnector[13] = fifoOut[48][0];
              muxOutConnector[14] = fifoOut[49][0];
              muxOutConnector[15] = fifoOut[50][0];
              muxOutConnector[16] = fifoOut[51][0];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       14: begin
              muxOutConnector[0] = fifoOut[35][0];
              muxOutConnector[1] = fifoOut[36][0];
              muxOutConnector[2] = fifoOut[37][0];
              muxOutConnector[3] = fifoOut[38][0];
              muxOutConnector[4] = fifoOut[39][0];
              muxOutConnector[5] = fifoOut[40][0];
              muxOutConnector[6] = fifoOut[41][0];
              muxOutConnector[7] = fifoOut[42][0];
              muxOutConnector[8] = fifoOut[43][0];
              muxOutConnector[9] = fifoOut[44][0];
              muxOutConnector[10] = fifoOut[45][0];
              muxOutConnector[11] = fifoOut[46][0];
              muxOutConnector[12] = fifoOut[47][0];
              muxOutConnector[13] = fifoOut[48][0];
              muxOutConnector[14] = fifoOut[49][0];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       15: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[2][13];
              muxOutConnector[18] = fifoOut[3][13];
              muxOutConnector[19] = fifoOut[4][13];
              muxOutConnector[20] = fifoOut[5][13];
              muxOutConnector[21] = fifoOut[6][13];
              muxOutConnector[22] = fifoOut[7][13];
              muxOutConnector[23] = fifoOut[8][13];
              muxOutConnector[24] = fifoOut[9][13];
              muxOutConnector[25] = fifoOut[10][13];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       16: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[2][13];
              muxOutConnector[18] = fifoOut[3][13];
              muxOutConnector[19] = fifoOut[4][13];
              muxOutConnector[20] = fifoOut[5][13];
              muxOutConnector[21] = fifoOut[6][13];
              muxOutConnector[22] = fifoOut[7][13];
              muxOutConnector[23] = fifoOut[8][13];
              muxOutConnector[24] = fifoOut[9][13];
              muxOutConnector[25] = fifoOut[10][13];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       17: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[2][13];
              muxOutConnector[18] = fifoOut[3][13];
              muxOutConnector[19] = fifoOut[4][13];
              muxOutConnector[20] = fifoOut[5][13];
              muxOutConnector[21] = fifoOut[6][13];
              muxOutConnector[22] = fifoOut[7][13];
              muxOutConnector[23] = fifoOut[8][13];
              muxOutConnector[24] = fifoOut[9][13];
              muxOutConnector[25] = fifoOut[10][13];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       18: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[2][13];
              muxOutConnector[18] = fifoOut[3][13];
              muxOutConnector[19] = fifoOut[4][13];
              muxOutConnector[20] = fifoOut[5][13];
              muxOutConnector[21] = fifoOut[6][13];
              muxOutConnector[22] = fifoOut[7][13];
              muxOutConnector[23] = fifoOut[8][13];
              muxOutConnector[24] = fifoOut[9][13];
              muxOutConnector[25] = fifoOut[10][13];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       19: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
