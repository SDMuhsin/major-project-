`timescale 1ns / 1ps
module LMem0To1_511_circ13_ys_scripted(
        muxOut,
        ly0In,
        wr_en,
        feedback_en,
        rd_address,
        rd_en,
        clk,
        rst
);
input feedback_en;
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 11;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        if(feedback_en) begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= fifoOut[i][c-1];
         end
        end
        else begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= ly0InConnector[i];
         end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[28][3];
              muxOutConnector[1] = fifoOut[29][3];
              muxOutConnector[2] = fifoOut[30][3];
              muxOutConnector[3] = fifoOut[31][3];
              muxOutConnector[4] = fifoOut[32][3];
              muxOutConnector[5] = fifoOut[33][3];
              muxOutConnector[6] = fifoOut[34][3];
              muxOutConnector[7] = fifoOut[35][3];
              muxOutConnector[8] = fifoOut[36][3];
              muxOutConnector[9] = fifoOut[37][3];
              muxOutConnector[10] = fifoOut[38][3];
              muxOutConnector[11] = fifoOut[39][3];
              muxOutConnector[12] = fifoOut[40][3];
              muxOutConnector[13] = fifoOut[41][3];
              muxOutConnector[14] = fifoOut[42][3];
              muxOutConnector[15] = fifoOut[43][3];
              muxOutConnector[16] = fifoOut[44][3];
              muxOutConnector[17] = fifoOut[45][3];
              muxOutConnector[18] = fifoOut[46][3];
              muxOutConnector[19] = fifoOut[47][3];
              muxOutConnector[20] = fifoOut[48][3];
              muxOutConnector[21] = fifoOut[49][3];
              muxOutConnector[22] = fifoOut[50][3];
              muxOutConnector[23] = fifoOut[51][3];
              muxOutConnector[24] = fifoOut[26][2];
              muxOutConnector[25] = fifoOut[27][2];
              muxOutConnector[26] = fifoOut[8][9];
              muxOutConnector[27] = fifoOut[9][9];
              muxOutConnector[28] = fifoOut[10][9];
              muxOutConnector[29] = fifoOut[11][9];
              muxOutConnector[30] = fifoOut[12][9];
              muxOutConnector[31] = fifoOut[13][9];
              muxOutConnector[32] = fifoOut[14][9];
              muxOutConnector[33] = fifoOut[15][9];
              muxOutConnector[34] = fifoOut[16][9];
              muxOutConnector[35] = fifoOut[17][9];
              muxOutConnector[36] = fifoOut[18][9];
              muxOutConnector[37] = fifoOut[19][9];
              muxOutConnector[38] = fifoOut[20][9];
              muxOutConnector[39] = fifoOut[21][9];
              muxOutConnector[40] = fifoOut[22][9];
              muxOutConnector[41] = fifoOut[23][9];
              muxOutConnector[42] = fifoOut[24][9];
              muxOutConnector[43] = fifoOut[25][9];
              muxOutConnector[44] = fifoOut[0][8];
              muxOutConnector[45] = fifoOut[1][8];
              muxOutConnector[46] = fifoOut[2][8];
              muxOutConnector[47] = fifoOut[3][8];
              muxOutConnector[48] = fifoOut[4][8];
              muxOutConnector[49] = fifoOut[5][8];
              muxOutConnector[50] = fifoOut[6][8];
              muxOutConnector[51] = fifoOut[7][8];
       end
       1: begin
              muxOutConnector[0] = fifoOut[28][3];
              muxOutConnector[1] = fifoOut[29][3];
              muxOutConnector[2] = fifoOut[30][3];
              muxOutConnector[3] = fifoOut[31][3];
              muxOutConnector[4] = fifoOut[32][3];
              muxOutConnector[5] = fifoOut[33][3];
              muxOutConnector[6] = fifoOut[34][3];
              muxOutConnector[7] = fifoOut[35][3];
              muxOutConnector[8] = fifoOut[36][3];
              muxOutConnector[9] = fifoOut[37][3];
              muxOutConnector[10] = fifoOut[38][3];
              muxOutConnector[11] = fifoOut[39][3];
              muxOutConnector[12] = fifoOut[40][3];
              muxOutConnector[13] = fifoOut[41][3];
              muxOutConnector[14] = fifoOut[42][3];
              muxOutConnector[15] = fifoOut[43][3];
              muxOutConnector[16] = fifoOut[44][3];
              muxOutConnector[17] = fifoOut[45][3];
              muxOutConnector[18] = fifoOut[46][3];
              muxOutConnector[19] = fifoOut[47][3];
              muxOutConnector[20] = fifoOut[48][3];
              muxOutConnector[21] = fifoOut[49][3];
              muxOutConnector[22] = fifoOut[50][3];
              muxOutConnector[23] = fifoOut[51][3];
              muxOutConnector[24] = fifoOut[26][2];
              muxOutConnector[25] = fifoOut[27][2];
              muxOutConnector[26] = fifoOut[8][9];
              muxOutConnector[27] = fifoOut[9][9];
              muxOutConnector[28] = fifoOut[10][9];
              muxOutConnector[29] = fifoOut[11][9];
              muxOutConnector[30] = fifoOut[12][9];
              muxOutConnector[31] = fifoOut[13][9];
              muxOutConnector[32] = fifoOut[14][9];
              muxOutConnector[33] = fifoOut[15][9];
              muxOutConnector[34] = fifoOut[16][9];
              muxOutConnector[35] = fifoOut[17][9];
              muxOutConnector[36] = fifoOut[18][9];
              muxOutConnector[37] = fifoOut[19][9];
              muxOutConnector[38] = fifoOut[20][9];
              muxOutConnector[39] = fifoOut[21][9];
              muxOutConnector[40] = fifoOut[22][9];
              muxOutConnector[41] = fifoOut[23][9];
              muxOutConnector[42] = fifoOut[24][9];
              muxOutConnector[43] = fifoOut[25][9];
              muxOutConnector[44] = fifoOut[0][8];
              muxOutConnector[45] = fifoOut[1][8];
              muxOutConnector[46] = fifoOut[2][8];
              muxOutConnector[47] = fifoOut[3][8];
              muxOutConnector[48] = fifoOut[4][8];
              muxOutConnector[49] = fifoOut[5][8];
              muxOutConnector[50] = fifoOut[6][8];
              muxOutConnector[51] = fifoOut[7][8];
       end
       2: begin
              muxOutConnector[0] = fifoOut[28][3];
              muxOutConnector[1] = fifoOut[29][3];
              muxOutConnector[2] = fifoOut[30][3];
              muxOutConnector[3] = fifoOut[31][3];
              muxOutConnector[4] = fifoOut[32][3];
              muxOutConnector[5] = fifoOut[33][3];
              muxOutConnector[6] = fifoOut[34][3];
              muxOutConnector[7] = fifoOut[35][3];
              muxOutConnector[8] = fifoOut[36][3];
              muxOutConnector[9] = fifoOut[37][3];
              muxOutConnector[10] = fifoOut[38][3];
              muxOutConnector[11] = fifoOut[39][3];
              muxOutConnector[12] = fifoOut[40][3];
              muxOutConnector[13] = fifoOut[41][3];
              muxOutConnector[14] = fifoOut[42][3];
              muxOutConnector[15] = fifoOut[43][3];
              muxOutConnector[16] = fifoOut[44][3];
              muxOutConnector[17] = fifoOut[45][3];
              muxOutConnector[18] = fifoOut[46][3];
              muxOutConnector[19] = fifoOut[47][3];
              muxOutConnector[20] = fifoOut[48][3];
              muxOutConnector[21] = fifoOut[49][3];
              muxOutConnector[22] = fifoOut[50][3];
              muxOutConnector[23] = fifoOut[51][3];
              muxOutConnector[24] = fifoOut[26][2];
              muxOutConnector[25] = fifoOut[27][2];
              muxOutConnector[26] = fifoOut[8][9];
              muxOutConnector[27] = fifoOut[9][9];
              muxOutConnector[28] = fifoOut[10][9];
              muxOutConnector[29] = fifoOut[11][9];
              muxOutConnector[30] = fifoOut[12][9];
              muxOutConnector[31] = fifoOut[13][9];
              muxOutConnector[32] = fifoOut[14][9];
              muxOutConnector[33] = fifoOut[15][9];
              muxOutConnector[34] = fifoOut[16][9];
              muxOutConnector[35] = fifoOut[17][9];
              muxOutConnector[36] = fifoOut[18][9];
              muxOutConnector[37] = fifoOut[19][9];
              muxOutConnector[38] = fifoOut[20][9];
              muxOutConnector[39] = fifoOut[21][9];
              muxOutConnector[40] = fifoOut[22][9];
              muxOutConnector[41] = fifoOut[23][9];
              muxOutConnector[42] = fifoOut[24][9];
              muxOutConnector[43] = fifoOut[25][9];
              muxOutConnector[44] = fifoOut[0][8];
              muxOutConnector[45] = fifoOut[1][8];
              muxOutConnector[46] = fifoOut[2][8];
              muxOutConnector[47] = fifoOut[3][8];
              muxOutConnector[48] = fifoOut[4][8];
              muxOutConnector[49] = fifoOut[5][8];
              muxOutConnector[50] = fifoOut[6][8];
              muxOutConnector[51] = fifoOut[7][8];
       end
       3: begin
              muxOutConnector[0] = fifoOut[28][3];
              muxOutConnector[1] = fifoOut[29][3];
              muxOutConnector[2] = fifoOut[30][3];
              muxOutConnector[3] = fifoOut[31][3];
              muxOutConnector[4] = fifoOut[32][3];
              muxOutConnector[5] = fifoOut[33][3];
              muxOutConnector[6] = fifoOut[34][3];
              muxOutConnector[7] = fifoOut[35][3];
              muxOutConnector[8] = fifoOut[36][3];
              muxOutConnector[9] = fifoOut[37][3];
              muxOutConnector[10] = fifoOut[38][3];
              muxOutConnector[11] = fifoOut[39][3];
              muxOutConnector[12] = fifoOut[40][3];
              muxOutConnector[13] = fifoOut[41][3];
              muxOutConnector[14] = fifoOut[42][3];
              muxOutConnector[15] = fifoOut[21][2];
              muxOutConnector[16] = fifoOut[22][2];
              muxOutConnector[17] = fifoOut[23][2];
              muxOutConnector[18] = fifoOut[24][2];
              muxOutConnector[19] = fifoOut[25][2];
              muxOutConnector[20] = fifoOut[0][1];
              muxOutConnector[21] = fifoOut[1][1];
              muxOutConnector[22] = fifoOut[2][1];
              muxOutConnector[23] = fifoOut[3][1];
              muxOutConnector[24] = fifoOut[4][1];
              muxOutConnector[25] = fifoOut[5][1];
              muxOutConnector[26] = fifoOut[8][9];
              muxOutConnector[27] = fifoOut[9][9];
              muxOutConnector[28] = fifoOut[10][9];
              muxOutConnector[29] = fifoOut[11][9];
              muxOutConnector[30] = fifoOut[12][9];
              muxOutConnector[31] = fifoOut[13][9];
              muxOutConnector[32] = fifoOut[14][9];
              muxOutConnector[33] = fifoOut[15][9];
              muxOutConnector[34] = fifoOut[16][9];
              muxOutConnector[35] = fifoOut[17][9];
              muxOutConnector[36] = fifoOut[18][9];
              muxOutConnector[37] = fifoOut[19][9];
              muxOutConnector[38] = fifoOut[20][9];
              muxOutConnector[39] = fifoOut[21][9];
              muxOutConnector[40] = fifoOut[22][9];
              muxOutConnector[41] = fifoOut[23][9];
              muxOutConnector[42] = fifoOut[24][9];
              muxOutConnector[43] = fifoOut[25][9];
              muxOutConnector[44] = fifoOut[0][8];
              muxOutConnector[45] = fifoOut[1][8];
              muxOutConnector[46] = fifoOut[2][8];
              muxOutConnector[47] = fifoOut[3][8];
              muxOutConnector[48] = fifoOut[4][8];
              muxOutConnector[49] = fifoOut[5][8];
              muxOutConnector[50] = fifoOut[6][8];
              muxOutConnector[51] = fifoOut[7][8];
       end
       4: begin
              muxOutConnector[0] = fifoOut[6][2];
              muxOutConnector[1] = fifoOut[7][2];
              muxOutConnector[2] = fifoOut[8][2];
              muxOutConnector[3] = fifoOut[9][2];
              muxOutConnector[4] = fifoOut[10][2];
              muxOutConnector[5] = fifoOut[11][2];
              muxOutConnector[6] = fifoOut[12][2];
              muxOutConnector[7] = fifoOut[13][2];
              muxOutConnector[8] = fifoOut[14][2];
              muxOutConnector[9] = fifoOut[15][2];
              muxOutConnector[10] = fifoOut[16][2];
              muxOutConnector[11] = fifoOut[17][2];
              muxOutConnector[12] = fifoOut[18][2];
              muxOutConnector[13] = fifoOut[19][2];
              muxOutConnector[14] = fifoOut[20][2];
              muxOutConnector[15] = fifoOut[21][2];
              muxOutConnector[16] = fifoOut[22][2];
              muxOutConnector[17] = fifoOut[23][2];
              muxOutConnector[18] = fifoOut[24][2];
              muxOutConnector[19] = fifoOut[25][2];
              muxOutConnector[20] = fifoOut[0][1];
              muxOutConnector[21] = fifoOut[1][1];
              muxOutConnector[22] = fifoOut[2][1];
              muxOutConnector[23] = fifoOut[3][1];
              muxOutConnector[24] = fifoOut[4][1];
              muxOutConnector[25] = fifoOut[5][1];
              muxOutConnector[26] = fifoOut[8][9];
              muxOutConnector[27] = fifoOut[9][9];
              muxOutConnector[28] = fifoOut[10][9];
              muxOutConnector[29] = fifoOut[11][9];
              muxOutConnector[30] = fifoOut[12][9];
              muxOutConnector[31] = fifoOut[13][9];
              muxOutConnector[32] = fifoOut[14][9];
              muxOutConnector[33] = fifoOut[15][9];
              muxOutConnector[34] = fifoOut[16][9];
              muxOutConnector[35] = fifoOut[17][9];
              muxOutConnector[36] = fifoOut[18][9];
              muxOutConnector[37] = fifoOut[19][9];
              muxOutConnector[38] = fifoOut[20][9];
              muxOutConnector[39] = fifoOut[21][9];
              muxOutConnector[40] = fifoOut[22][9];
              muxOutConnector[41] = fifoOut[23][9];
              muxOutConnector[42] = fifoOut[24][9];
              muxOutConnector[43] = fifoOut[25][9];
              muxOutConnector[44] = fifoOut[0][8];
              muxOutConnector[45] = fifoOut[1][8];
              muxOutConnector[46] = fifoOut[2][8];
              muxOutConnector[47] = fifoOut[3][8];
              muxOutConnector[48] = fifoOut[4][8];
              muxOutConnector[49] = fifoOut[5][8];
              muxOutConnector[50] = fifoOut[6][8];
              muxOutConnector[51] = fifoOut[7][8];
       end
       5: begin
              muxOutConnector[0] = fifoOut[6][2];
              muxOutConnector[1] = fifoOut[7][2];
              muxOutConnector[2] = fifoOut[8][2];
              muxOutConnector[3] = fifoOut[9][2];
              muxOutConnector[4] = fifoOut[10][2];
              muxOutConnector[5] = fifoOut[11][2];
              muxOutConnector[6] = fifoOut[12][2];
              muxOutConnector[7] = fifoOut[13][2];
              muxOutConnector[8] = fifoOut[14][2];
              muxOutConnector[9] = fifoOut[15][2];
              muxOutConnector[10] = fifoOut[16][2];
              muxOutConnector[11] = fifoOut[17][2];
              muxOutConnector[12] = fifoOut[18][2];
              muxOutConnector[13] = fifoOut[19][2];
              muxOutConnector[14] = fifoOut[20][2];
              muxOutConnector[15] = fifoOut[21][2];
              muxOutConnector[16] = fifoOut[22][2];
              muxOutConnector[17] = fifoOut[23][2];
              muxOutConnector[18] = fifoOut[24][2];
              muxOutConnector[19] = fifoOut[25][2];
              muxOutConnector[20] = fifoOut[0][1];
              muxOutConnector[21] = fifoOut[1][1];
              muxOutConnector[22] = fifoOut[2][1];
              muxOutConnector[23] = fifoOut[3][1];
              muxOutConnector[24] = fifoOut[4][1];
              muxOutConnector[25] = fifoOut[5][1];
              muxOutConnector[26] = fifoOut[8][9];
              muxOutConnector[27] = fifoOut[9][9];
              muxOutConnector[28] = fifoOut[10][9];
              muxOutConnector[29] = fifoOut[11][9];
              muxOutConnector[30] = fifoOut[12][9];
              muxOutConnector[31] = fifoOut[13][9];
              muxOutConnector[32] = fifoOut[14][9];
              muxOutConnector[33] = fifoOut[15][9];
              muxOutConnector[34] = fifoOut[16][9];
              muxOutConnector[35] = fifoOut[17][9];
              muxOutConnector[36] = fifoOut[18][9];
              muxOutConnector[37] = fifoOut[19][9];
              muxOutConnector[38] = fifoOut[20][9];
              muxOutConnector[39] = fifoOut[21][9];
              muxOutConnector[40] = fifoOut[22][9];
              muxOutConnector[41] = fifoOut[23][9];
              muxOutConnector[42] = fifoOut[24][9];
              muxOutConnector[43] = fifoOut[25][9];
              muxOutConnector[44] = fifoOut[0][8];
              muxOutConnector[45] = fifoOut[1][8];
              muxOutConnector[46] = fifoOut[2][8];
              muxOutConnector[47] = fifoOut[3][8];
              muxOutConnector[48] = fifoOut[4][8];
              muxOutConnector[49] = fifoOut[5][8];
              muxOutConnector[50] = fifoOut[6][8];
              muxOutConnector[51] = fifoOut[7][8];
       end
       6: begin
              muxOutConnector[0] = fifoOut[6][2];
              muxOutConnector[1] = fifoOut[7][2];
              muxOutConnector[2] = fifoOut[8][2];
              muxOutConnector[3] = fifoOut[9][2];
              muxOutConnector[4] = fifoOut[10][2];
              muxOutConnector[5] = fifoOut[11][2];
              muxOutConnector[6] = fifoOut[12][2];
              muxOutConnector[7] = fifoOut[13][2];
              muxOutConnector[8] = fifoOut[14][2];
              muxOutConnector[9] = fifoOut[15][2];
              muxOutConnector[10] = fifoOut[16][2];
              muxOutConnector[11] = fifoOut[17][2];
              muxOutConnector[12] = fifoOut[18][2];
              muxOutConnector[13] = fifoOut[19][2];
              muxOutConnector[14] = fifoOut[20][2];
              muxOutConnector[15] = fifoOut[21][2];
              muxOutConnector[16] = fifoOut[22][2];
              muxOutConnector[17] = fifoOut[23][2];
              muxOutConnector[18] = fifoOut[24][2];
              muxOutConnector[19] = fifoOut[25][2];
              muxOutConnector[20] = fifoOut[0][1];
              muxOutConnector[21] = fifoOut[1][1];
              muxOutConnector[22] = fifoOut[2][1];
              muxOutConnector[23] = fifoOut[3][1];
              muxOutConnector[24] = fifoOut[4][1];
              muxOutConnector[25] = fifoOut[5][1];
              muxOutConnector[26] = fifoOut[8][9];
              muxOutConnector[27] = fifoOut[9][9];
              muxOutConnector[28] = fifoOut[10][9];
              muxOutConnector[29] = fifoOut[11][9];
              muxOutConnector[30] = fifoOut[12][9];
              muxOutConnector[31] = fifoOut[13][9];
              muxOutConnector[32] = fifoOut[14][9];
              muxOutConnector[33] = fifoOut[15][9];
              muxOutConnector[34] = fifoOut[16][9];
              muxOutConnector[35] = fifoOut[17][9];
              muxOutConnector[36] = fifoOut[18][9];
              muxOutConnector[37] = fifoOut[19][9];
              muxOutConnector[38] = fifoOut[20][9];
              muxOutConnector[39] = fifoOut[21][9];
              muxOutConnector[40] = fifoOut[22][9];
              muxOutConnector[41] = fifoOut[23][9];
              muxOutConnector[42] = fifoOut[24][9];
              muxOutConnector[43] = fifoOut[25][9];
              muxOutConnector[44] = fifoOut[0][8];
              muxOutConnector[45] = fifoOut[1][8];
              muxOutConnector[46] = fifoOut[2][8];
              muxOutConnector[47] = fifoOut[3][8];
              muxOutConnector[48] = fifoOut[4][8];
              muxOutConnector[49] = fifoOut[5][8];
              muxOutConnector[50] = fifoOut[6][8];
              muxOutConnector[51] = fifoOut[7][8];
       end
       7: begin
              muxOutConnector[0] = fifoOut[6][2];
              muxOutConnector[1] = fifoOut[7][2];
              muxOutConnector[2] = fifoOut[8][2];
              muxOutConnector[3] = fifoOut[9][2];
              muxOutConnector[4] = fifoOut[10][2];
              muxOutConnector[5] = fifoOut[11][2];
              muxOutConnector[6] = fifoOut[12][2];
              muxOutConnector[7] = fifoOut[13][2];
              muxOutConnector[8] = fifoOut[14][2];
              muxOutConnector[9] = fifoOut[15][2];
              muxOutConnector[10] = fifoOut[16][2];
              muxOutConnector[11] = fifoOut[17][2];
              muxOutConnector[12] = fifoOut[18][2];
              muxOutConnector[13] = fifoOut[19][2];
              muxOutConnector[14] = fifoOut[20][2];
              muxOutConnector[15] = fifoOut[21][2];
              muxOutConnector[16] = fifoOut[22][2];
              muxOutConnector[17] = fifoOut[23][2];
              muxOutConnector[18] = fifoOut[24][2];
              muxOutConnector[19] = fifoOut[25][2];
              muxOutConnector[20] = fifoOut[0][1];
              muxOutConnector[21] = fifoOut[1][1];
              muxOutConnector[22] = fifoOut[2][1];
              muxOutConnector[23] = fifoOut[3][1];
              muxOutConnector[24] = fifoOut[4][1];
              muxOutConnector[25] = fifoOut[5][1];
              muxOutConnector[26] = fifoOut[8][9];
              muxOutConnector[27] = fifoOut[9][9];
              muxOutConnector[28] = fifoOut[10][9];
              muxOutConnector[29] = fifoOut[11][9];
              muxOutConnector[30] = fifoOut[12][9];
              muxOutConnector[31] = fifoOut[13][9];
              muxOutConnector[32] = fifoOut[14][9];
              muxOutConnector[33] = fifoOut[15][9];
              muxOutConnector[34] = fifoOut[16][9];
              muxOutConnector[35] = fifoOut[17][9];
              muxOutConnector[36] = fifoOut[18][9];
              muxOutConnector[37] = fifoOut[19][9];
              muxOutConnector[38] = fifoOut[20][9];
              muxOutConnector[39] = fifoOut[21][9];
              muxOutConnector[40] = fifoOut[22][9];
              muxOutConnector[41] = fifoOut[23][9];
              muxOutConnector[42] = fifoOut[24][9];
              muxOutConnector[43] = fifoOut[25][9];
              muxOutConnector[44] = fifoOut[0][8];
              muxOutConnector[45] = fifoOut[1][8];
              muxOutConnector[46] = fifoOut[2][8];
              muxOutConnector[47] = fifoOut[3][8];
              muxOutConnector[48] = fifoOut[4][8];
              muxOutConnector[49] = fifoOut[5][8];
              muxOutConnector[50] = fifoOut[6][8];
              muxOutConnector[51] = fifoOut[7][8];
       end
       8: begin
              muxOutConnector[0] = fifoOut[6][2];
              muxOutConnector[1] = fifoOut[7][2];
              muxOutConnector[2] = fifoOut[8][2];
              muxOutConnector[3] = fifoOut[9][2];
              muxOutConnector[4] = fifoOut[10][2];
              muxOutConnector[5] = fifoOut[11][2];
              muxOutConnector[6] = fifoOut[12][2];
              muxOutConnector[7] = fifoOut[13][2];
              muxOutConnector[8] = fifoOut[14][2];
              muxOutConnector[9] = fifoOut[15][2];
              muxOutConnector[10] = fifoOut[16][2];
              muxOutConnector[11] = fifoOut[17][2];
              muxOutConnector[12] = fifoOut[18][2];
              muxOutConnector[13] = fifoOut[19][2];
              muxOutConnector[14] = fifoOut[20][2];
              muxOutConnector[15] = fifoOut[21][2];
              muxOutConnector[16] = fifoOut[22][2];
              muxOutConnector[17] = fifoOut[23][2];
              muxOutConnector[18] = fifoOut[24][2];
              muxOutConnector[19] = fifoOut[25][2];
              muxOutConnector[20] = fifoOut[0][1];
              muxOutConnector[21] = fifoOut[1][1];
              muxOutConnector[22] = fifoOut[2][1];
              muxOutConnector[23] = fifoOut[3][1];
              muxOutConnector[24] = fifoOut[4][1];
              muxOutConnector[25] = fifoOut[5][1];
              muxOutConnector[26] = fifoOut[8][9];
              muxOutConnector[27] = fifoOut[9][9];
              muxOutConnector[28] = fifoOut[10][9];
              muxOutConnector[29] = fifoOut[11][9];
              muxOutConnector[30] = fifoOut[12][9];
              muxOutConnector[31] = fifoOut[13][9];
              muxOutConnector[32] = fifoOut[14][9];
              muxOutConnector[33] = fifoOut[15][9];
              muxOutConnector[34] = fifoOut[16][9];
              muxOutConnector[35] = fifoOut[17][9];
              muxOutConnector[36] = fifoOut[18][9];
              muxOutConnector[37] = fifoOut[19][9];
              muxOutConnector[38] = fifoOut[20][9];
              muxOutConnector[39] = fifoOut[21][9];
              muxOutConnector[40] = fifoOut[22][9];
              muxOutConnector[41] = fifoOut[23][9];
              muxOutConnector[42] = fifoOut[24][9];
              muxOutConnector[43] = fifoOut[25][9];
              muxOutConnector[44] = fifoOut[0][8];
              muxOutConnector[45] = fifoOut[1][8];
              muxOutConnector[46] = fifoOut[2][8];
              muxOutConnector[47] = fifoOut[3][8];
              muxOutConnector[48] = fifoOut[4][8];
              muxOutConnector[49] = fifoOut[5][8];
              muxOutConnector[50] = fifoOut[6][8];
              muxOutConnector[51] = fifoOut[7][8];
       end
       9: begin
              muxOutConnector[0] = fifoOut[6][2];
              muxOutConnector[1] = fifoOut[7][2];
              muxOutConnector[2] = fifoOut[8][2];
              muxOutConnector[3] = fifoOut[9][2];
              muxOutConnector[4] = fifoOut[10][2];
              muxOutConnector[5] = fifoOut[11][2];
              muxOutConnector[6] = fifoOut[12][2];
              muxOutConnector[7] = fifoOut[13][2];
              muxOutConnector[8] = fifoOut[14][2];
              muxOutConnector[9] = fifoOut[15][2];
              muxOutConnector[10] = fifoOut[16][2];
              muxOutConnector[11] = fifoOut[17][2];
              muxOutConnector[12] = fifoOut[18][2];
              muxOutConnector[13] = fifoOut[19][2];
              muxOutConnector[14] = fifoOut[20][2];
              muxOutConnector[15] = fifoOut[21][2];
              muxOutConnector[16] = fifoOut[22][2];
              muxOutConnector[17] = fifoOut[23][2];
              muxOutConnector[18] = fifoOut[24][2];
              muxOutConnector[19] = fifoOut[25][2];
              muxOutConnector[20] = fifoOut[0][1];
              muxOutConnector[21] = fifoOut[1][1];
              muxOutConnector[22] = fifoOut[2][1];
              muxOutConnector[23] = fifoOut[3][1];
              muxOutConnector[24] = fifoOut[4][1];
              muxOutConnector[25] = fifoOut[5][1];
              muxOutConnector[26] = fifoOut[8][9];
              muxOutConnector[27] = fifoOut[9][9];
              muxOutConnector[28] = fifoOut[10][9];
              muxOutConnector[29] = fifoOut[11][9];
              muxOutConnector[30] = fifoOut[12][9];
              muxOutConnector[31] = fifoOut[13][9];
              muxOutConnector[32] = fifoOut[14][9];
              muxOutConnector[33] = fifoOut[15][9];
              muxOutConnector[34] = fifoOut[16][9];
              muxOutConnector[35] = fifoOut[48][8];
              muxOutConnector[36] = fifoOut[49][8];
              muxOutConnector[37] = fifoOut[50][8];
              muxOutConnector[38] = fifoOut[51][8];
              muxOutConnector[39] = fifoOut[26][7];
              muxOutConnector[40] = fifoOut[27][7];
              muxOutConnector[41] = fifoOut[28][7];
              muxOutConnector[42] = fifoOut[29][7];
              muxOutConnector[43] = fifoOut[30][7];
              muxOutConnector[44] = fifoOut[31][7];
              muxOutConnector[45] = fifoOut[32][7];
              muxOutConnector[46] = fifoOut[33][7];
              muxOutConnector[47] = fifoOut[34][7];
              muxOutConnector[48] = fifoOut[35][7];
              muxOutConnector[49] = fifoOut[36][7];
              muxOutConnector[50] = fifoOut[37][7];
              muxOutConnector[51] = fifoOut[38][7];
       end
       10: begin
              muxOutConnector[0] = fifoOut[6][2];
              muxOutConnector[1] = fifoOut[7][2];
              muxOutConnector[2] = fifoOut[8][2];
              muxOutConnector[3] = fifoOut[9][2];
              muxOutConnector[4] = fifoOut[10][2];
              muxOutConnector[5] = fifoOut[11][2];
              muxOutConnector[6] = fifoOut[12][2];
              muxOutConnector[7] = fifoOut[13][2];
              muxOutConnector[8] = fifoOut[14][2];
              muxOutConnector[9] = fifoOut[15][2];
              muxOutConnector[10] = fifoOut[16][2];
              muxOutConnector[11] = fifoOut[17][2];
              muxOutConnector[12] = fifoOut[18][2];
              muxOutConnector[13] = fifoOut[19][2];
              muxOutConnector[14] = fifoOut[20][2];
              muxOutConnector[15] = fifoOut[21][2];
              muxOutConnector[16] = fifoOut[22][2];
              muxOutConnector[17] = fifoOut[23][2];
              muxOutConnector[18] = fifoOut[24][2];
              muxOutConnector[19] = fifoOut[25][2];
              muxOutConnector[20] = fifoOut[0][1];
              muxOutConnector[21] = fifoOut[1][1];
              muxOutConnector[22] = fifoOut[2][1];
              muxOutConnector[23] = fifoOut[3][1];
              muxOutConnector[24] = fifoOut[4][1];
              muxOutConnector[25] = fifoOut[5][1];
              muxOutConnector[26] = fifoOut[39][8];
              muxOutConnector[27] = fifoOut[40][8];
              muxOutConnector[28] = fifoOut[41][8];
              muxOutConnector[29] = fifoOut[42][8];
              muxOutConnector[30] = fifoOut[43][8];
              muxOutConnector[31] = fifoOut[44][8];
              muxOutConnector[32] = fifoOut[45][8];
              muxOutConnector[33] = fifoOut[46][8];
              muxOutConnector[34] = fifoOut[47][8];
              muxOutConnector[35] = fifoOut[48][8];
              muxOutConnector[36] = fifoOut[49][8];
              muxOutConnector[37] = fifoOut[50][8];
              muxOutConnector[38] = fifoOut[51][8];
              muxOutConnector[39] = fifoOut[26][7];
              muxOutConnector[40] = fifoOut[27][7];
              muxOutConnector[41] = fifoOut[28][7];
              muxOutConnector[42] = fifoOut[29][7];
              muxOutConnector[43] = fifoOut[30][7];
              muxOutConnector[44] = fifoOut[31][7];
              muxOutConnector[45] = fifoOut[32][7];
              muxOutConnector[46] = fifoOut[33][7];
              muxOutConnector[47] = fifoOut[34][7];
              muxOutConnector[48] = fifoOut[35][7];
              muxOutConnector[49] = fifoOut[36][7];
              muxOutConnector[50] = fifoOut[37][7];
              muxOutConnector[51] = fifoOut[38][7];
       end
       11: begin
              muxOutConnector[0] = fifoOut[6][2];
              muxOutConnector[1] = fifoOut[7][2];
              muxOutConnector[2] = fifoOut[8][2];
              muxOutConnector[3] = fifoOut[9][2];
              muxOutConnector[4] = fifoOut[10][2];
              muxOutConnector[5] = fifoOut[11][2];
              muxOutConnector[6] = fifoOut[12][2];
              muxOutConnector[7] = fifoOut[13][2];
              muxOutConnector[8] = fifoOut[14][2];
              muxOutConnector[9] = fifoOut[15][2];
              muxOutConnector[10] = fifoOut[16][2];
              muxOutConnector[11] = fifoOut[17][2];
              muxOutConnector[12] = fifoOut[18][2];
              muxOutConnector[13] = fifoOut[19][2];
              muxOutConnector[14] = fifoOut[20][2];
              muxOutConnector[15] = fifoOut[21][2];
              muxOutConnector[16] = fifoOut[22][2];
              muxOutConnector[17] = fifoOut[23][2];
              muxOutConnector[18] = fifoOut[24][2];
              muxOutConnector[19] = fifoOut[25][2];
              muxOutConnector[20] = fifoOut[0][1];
              muxOutConnector[21] = fifoOut[1][1];
              muxOutConnector[22] = fifoOut[2][1];
              muxOutConnector[23] = fifoOut[3][1];
              muxOutConnector[24] = fifoOut[4][1];
              muxOutConnector[25] = fifoOut[5][1];
              muxOutConnector[26] = fifoOut[39][8];
              muxOutConnector[27] = fifoOut[40][8];
              muxOutConnector[28] = fifoOut[41][8];
              muxOutConnector[29] = fifoOut[42][8];
              muxOutConnector[30] = fifoOut[43][8];
              muxOutConnector[31] = fifoOut[44][8];
              muxOutConnector[32] = fifoOut[45][8];
              muxOutConnector[33] = fifoOut[46][8];
              muxOutConnector[34] = fifoOut[47][8];
              muxOutConnector[35] = fifoOut[48][8];
              muxOutConnector[36] = fifoOut[49][8];
              muxOutConnector[37] = fifoOut[50][8];
              muxOutConnector[38] = fifoOut[51][8];
              muxOutConnector[39] = fifoOut[26][7];
              muxOutConnector[40] = fifoOut[27][7];
              muxOutConnector[41] = fifoOut[28][7];
              muxOutConnector[42] = fifoOut[29][7];
              muxOutConnector[43] = fifoOut[30][7];
              muxOutConnector[44] = fifoOut[31][7];
              muxOutConnector[45] = fifoOut[32][7];
              muxOutConnector[46] = fifoOut[33][7];
              muxOutConnector[47] = fifoOut[34][7];
              muxOutConnector[48] = fifoOut[35][7];
              muxOutConnector[49] = fifoOut[36][7];
              muxOutConnector[50] = fifoOut[37][7];
              muxOutConnector[51] = fifoOut[38][7];
       end
       12: begin
              muxOutConnector[0] = fifoOut[6][2];
              muxOutConnector[1] = fifoOut[7][2];
              muxOutConnector[2] = fifoOut[8][2];
              muxOutConnector[3] = fifoOut[9][2];
              muxOutConnector[4] = fifoOut[10][2];
              muxOutConnector[5] = fifoOut[11][2];
              muxOutConnector[6] = fifoOut[12][2];
              muxOutConnector[7] = fifoOut[13][2];
              muxOutConnector[8] = fifoOut[14][2];
              muxOutConnector[9] = fifoOut[15][2];
              muxOutConnector[10] = fifoOut[16][2];
              muxOutConnector[11] = fifoOut[17][2];
              muxOutConnector[12] = fifoOut[18][2];
              muxOutConnector[13] = fifoOut[19][2];
              muxOutConnector[14] = fifoOut[20][2];
              muxOutConnector[15] = fifoOut[21][2];
              muxOutConnector[16] = fifoOut[22][2];
              muxOutConnector[17] = fifoOut[23][2];
              muxOutConnector[18] = fifoOut[24][2];
              muxOutConnector[19] = fifoOut[25][2];
              muxOutConnector[20] = fifoOut[0][1];
              muxOutConnector[21] = fifoOut[1][1];
              muxOutConnector[22] = fifoOut[2][1];
              muxOutConnector[23] = fifoOut[3][1];
              muxOutConnector[24] = fifoOut[4][1];
              muxOutConnector[25] = fifoOut[5][1];
              muxOutConnector[26] = fifoOut[39][8];
              muxOutConnector[27] = fifoOut[40][8];
              muxOutConnector[28] = fifoOut[41][8];
              muxOutConnector[29] = fifoOut[42][8];
              muxOutConnector[30] = fifoOut[43][8];
              muxOutConnector[31] = fifoOut[44][8];
              muxOutConnector[32] = fifoOut[45][8];
              muxOutConnector[33] = fifoOut[46][8];
              muxOutConnector[34] = fifoOut[47][8];
              muxOutConnector[35] = fifoOut[48][8];
              muxOutConnector[36] = fifoOut[49][8];
              muxOutConnector[37] = fifoOut[50][8];
              muxOutConnector[38] = fifoOut[51][8];
              muxOutConnector[39] = fifoOut[26][7];
              muxOutConnector[40] = fifoOut[27][7];
              muxOutConnector[41] = fifoOut[28][7];
              muxOutConnector[42] = fifoOut[29][7];
              muxOutConnector[43] = fifoOut[30][7];
              muxOutConnector[44] = fifoOut[31][7];
              muxOutConnector[45] = fifoOut[32][7];
              muxOutConnector[46] = fifoOut[33][7];
              muxOutConnector[47] = fifoOut[34][7];
              muxOutConnector[48] = fifoOut[35][7];
              muxOutConnector[49] = fifoOut[36][7];
              muxOutConnector[50] = fifoOut[37][7];
              muxOutConnector[51] = fifoOut[38][7];
       end
       13: begin
              muxOutConnector[0] = fifoOut[6][2];
              muxOutConnector[1] = fifoOut[7][2];
              muxOutConnector[2] = fifoOut[8][2];
              muxOutConnector[3] = fifoOut[9][2];
              muxOutConnector[4] = fifoOut[10][2];
              muxOutConnector[5] = fifoOut[11][2];
              muxOutConnector[6] = fifoOut[12][2];
              muxOutConnector[7] = fifoOut[13][2];
              muxOutConnector[8] = fifoOut[14][2];
              muxOutConnector[9] = fifoOut[15][2];
              muxOutConnector[10] = fifoOut[16][2];
              muxOutConnector[11] = fifoOut[48][1];
              muxOutConnector[12] = fifoOut[49][1];
              muxOutConnector[13] = fifoOut[50][1];
              muxOutConnector[14] = fifoOut[51][1];
              muxOutConnector[15] = fifoOut[26][0];
              muxOutConnector[16] = fifoOut[27][0];
              muxOutConnector[17] = fifoOut[28][0];
              muxOutConnector[18] = fifoOut[29][0];
              muxOutConnector[19] = fifoOut[30][0];
              muxOutConnector[20] = fifoOut[31][0];
              muxOutConnector[21] = fifoOut[32][0];
              muxOutConnector[22] = fifoOut[33][0];
              muxOutConnector[23] = fifoOut[34][0];
              muxOutConnector[24] = fifoOut[35][0];
              muxOutConnector[25] = fifoOut[36][0];
              muxOutConnector[26] = fifoOut[39][8];
              muxOutConnector[27] = fifoOut[40][8];
              muxOutConnector[28] = fifoOut[41][8];
              muxOutConnector[29] = fifoOut[42][8];
              muxOutConnector[30] = fifoOut[43][8];
              muxOutConnector[31] = fifoOut[44][8];
              muxOutConnector[32] = fifoOut[45][8];
              muxOutConnector[33] = fifoOut[46][8];
              muxOutConnector[34] = fifoOut[47][8];
              muxOutConnector[35] = fifoOut[48][8];
              muxOutConnector[36] = fifoOut[49][8];
              muxOutConnector[37] = fifoOut[50][8];
              muxOutConnector[38] = fifoOut[51][8];
              muxOutConnector[39] = fifoOut[26][7];
              muxOutConnector[40] = fifoOut[27][7];
              muxOutConnector[41] = fifoOut[28][7];
              muxOutConnector[42] = fifoOut[29][7];
              muxOutConnector[43] = fifoOut[30][7];
              muxOutConnector[44] = fifoOut[31][7];
              muxOutConnector[45] = fifoOut[32][7];
              muxOutConnector[46] = fifoOut[33][7];
              muxOutConnector[47] = fifoOut[34][7];
              muxOutConnector[48] = fifoOut[35][7];
              muxOutConnector[49] = fifoOut[36][7];
              muxOutConnector[50] = fifoOut[37][7];
              muxOutConnector[51] = fifoOut[38][7];
       end
       14: begin
              muxOutConnector[0] = fifoOut[37][1];
              muxOutConnector[1] = fifoOut[38][1];
              muxOutConnector[2] = fifoOut[39][1];
              muxOutConnector[3] = fifoOut[40][1];
              muxOutConnector[4] = fifoOut[41][1];
              muxOutConnector[5] = fifoOut[42][1];
              muxOutConnector[6] = fifoOut[43][1];
              muxOutConnector[7] = fifoOut[44][1];
              muxOutConnector[8] = fifoOut[45][1];
              muxOutConnector[9] = fifoOut[46][1];
              muxOutConnector[10] = fifoOut[47][1];
              muxOutConnector[11] = fifoOut[48][1];
              muxOutConnector[12] = fifoOut[49][1];
              muxOutConnector[13] = fifoOut[50][1];
              muxOutConnector[14] = fifoOut[51][1];
              muxOutConnector[15] = fifoOut[26][0];
              muxOutConnector[16] = fifoOut[27][0];
              muxOutConnector[17] = fifoOut[28][0];
              muxOutConnector[18] = fifoOut[29][0];
              muxOutConnector[19] = fifoOut[30][0];
              muxOutConnector[20] = fifoOut[31][0];
              muxOutConnector[21] = fifoOut[32][0];
              muxOutConnector[22] = fifoOut[33][0];
              muxOutConnector[23] = fifoOut[34][0];
              muxOutConnector[24] = fifoOut[35][0];
              muxOutConnector[25] = fifoOut[36][0];
              muxOutConnector[26] = fifoOut[39][8];
              muxOutConnector[27] = fifoOut[40][8];
              muxOutConnector[28] = fifoOut[41][8];
              muxOutConnector[29] = fifoOut[42][8];
              muxOutConnector[30] = fifoOut[43][8];
              muxOutConnector[31] = fifoOut[44][8];
              muxOutConnector[32] = fifoOut[45][8];
              muxOutConnector[33] = fifoOut[46][8];
              muxOutConnector[34] = fifoOut[47][8];
              muxOutConnector[35] = fifoOut[48][8];
              muxOutConnector[36] = fifoOut[49][8];
              muxOutConnector[37] = fifoOut[50][8];
              muxOutConnector[38] = fifoOut[51][8];
              muxOutConnector[39] = fifoOut[26][7];
              muxOutConnector[40] = fifoOut[27][7];
              muxOutConnector[41] = fifoOut[28][7];
              muxOutConnector[42] = fifoOut[29][7];
              muxOutConnector[43] = fifoOut[30][7];
              muxOutConnector[44] = fifoOut[31][7];
              muxOutConnector[45] = fifoOut[32][7];
              muxOutConnector[46] = fifoOut[33][7];
              muxOutConnector[47] = fifoOut[34][7];
              muxOutConnector[48] = fifoOut[35][7];
              muxOutConnector[49] = fifoOut[36][7];
              muxOutConnector[50] = fifoOut[37][7];
              muxOutConnector[51] = fifoOut[38][7];
       end
       15: begin
              muxOutConnector[0] = fifoOut[37][1];
              muxOutConnector[1] = fifoOut[38][1];
              muxOutConnector[2] = fifoOut[39][1];
              muxOutConnector[3] = fifoOut[40][1];
              muxOutConnector[4] = fifoOut[41][1];
              muxOutConnector[5] = fifoOut[42][1];
              muxOutConnector[6] = fifoOut[43][1];
              muxOutConnector[7] = fifoOut[44][1];
              muxOutConnector[8] = fifoOut[45][1];
              muxOutConnector[9] = fifoOut[46][1];
              muxOutConnector[10] = fifoOut[47][1];
              muxOutConnector[11] = fifoOut[48][1];
              muxOutConnector[12] = fifoOut[49][1];
              muxOutConnector[13] = fifoOut[50][1];
              muxOutConnector[14] = fifoOut[51][1];
              muxOutConnector[15] = fifoOut[26][0];
              muxOutConnector[16] = fifoOut[27][0];
              muxOutConnector[17] = fifoOut[28][0];
              muxOutConnector[18] = fifoOut[29][0];
              muxOutConnector[19] = fifoOut[30][0];
              muxOutConnector[20] = fifoOut[31][0];
              muxOutConnector[21] = fifoOut[32][0];
              muxOutConnector[22] = fifoOut[33][0];
              muxOutConnector[23] = fifoOut[34][0];
              muxOutConnector[24] = fifoOut[35][0];
              muxOutConnector[25] = fifoOut[36][0];
              muxOutConnector[26] = fifoOut[39][8];
              muxOutConnector[27] = fifoOut[40][8];
              muxOutConnector[28] = fifoOut[41][8];
              muxOutConnector[29] = fifoOut[42][8];
              muxOutConnector[30] = fifoOut[43][8];
              muxOutConnector[31] = fifoOut[44][8];
              muxOutConnector[32] = fifoOut[45][8];
              muxOutConnector[33] = fifoOut[46][8];
              muxOutConnector[34] = fifoOut[47][8];
              muxOutConnector[35] = fifoOut[48][8];
              muxOutConnector[36] = fifoOut[49][8];
              muxOutConnector[37] = fifoOut[50][8];
              muxOutConnector[38] = fifoOut[51][8];
              muxOutConnector[39] = fifoOut[26][7];
              muxOutConnector[40] = fifoOut[27][7];
              muxOutConnector[41] = fifoOut[28][7];
              muxOutConnector[42] = fifoOut[29][7];
              muxOutConnector[43] = fifoOut[30][7];
              muxOutConnector[44] = fifoOut[31][7];
              muxOutConnector[45] = fifoOut[32][7];
              muxOutConnector[46] = fifoOut[33][7];
              muxOutConnector[47] = fifoOut[34][7];
              muxOutConnector[48] = fifoOut[35][7];
              muxOutConnector[49] = fifoOut[36][7];
              muxOutConnector[50] = fifoOut[37][7];
              muxOutConnector[51] = fifoOut[38][7];
       end
       16: begin
              muxOutConnector[0] = fifoOut[37][1];
              muxOutConnector[1] = fifoOut[38][1];
              muxOutConnector[2] = fifoOut[39][1];
              muxOutConnector[3] = fifoOut[40][1];
              muxOutConnector[4] = fifoOut[41][1];
              muxOutConnector[5] = fifoOut[42][1];
              muxOutConnector[6] = fifoOut[43][1];
              muxOutConnector[7] = fifoOut[44][1];
              muxOutConnector[8] = fifoOut[45][1];
              muxOutConnector[9] = fifoOut[46][1];
              muxOutConnector[10] = fifoOut[47][1];
              muxOutConnector[11] = fifoOut[48][1];
              muxOutConnector[12] = fifoOut[49][1];
              muxOutConnector[13] = fifoOut[50][1];
              muxOutConnector[14] = fifoOut[51][1];
              muxOutConnector[15] = fifoOut[26][0];
              muxOutConnector[16] = fifoOut[27][0];
              muxOutConnector[17] = fifoOut[28][0];
              muxOutConnector[18] = fifoOut[29][0];
              muxOutConnector[19] = fifoOut[30][0];
              muxOutConnector[20] = fifoOut[31][0];
              muxOutConnector[21] = fifoOut[32][0];
              muxOutConnector[22] = fifoOut[33][0];
              muxOutConnector[23] = fifoOut[34][0];
              muxOutConnector[24] = fifoOut[35][0];
              muxOutConnector[25] = fifoOut[36][0];
              muxOutConnector[26] = fifoOut[39][8];
              muxOutConnector[27] = fifoOut[40][8];
              muxOutConnector[28] = fifoOut[41][8];
              muxOutConnector[29] = fifoOut[42][8];
              muxOutConnector[30] = fifoOut[43][8];
              muxOutConnector[31] = fifoOut[44][8];
              muxOutConnector[32] = fifoOut[45][8];
              muxOutConnector[33] = fifoOut[46][8];
              muxOutConnector[34] = fifoOut[47][8];
              muxOutConnector[35] = fifoOut[48][8];
              muxOutConnector[36] = fifoOut[49][8];
              muxOutConnector[37] = fifoOut[50][8];
              muxOutConnector[38] = fifoOut[51][8];
              muxOutConnector[39] = fifoOut[26][7];
              muxOutConnector[40] = fifoOut[27][7];
              muxOutConnector[41] = fifoOut[28][7];
              muxOutConnector[42] = fifoOut[29][7];
              muxOutConnector[43] = fifoOut[30][7];
              muxOutConnector[44] = fifoOut[31][7];
              muxOutConnector[45] = fifoOut[32][7];
              muxOutConnector[46] = fifoOut[33][7];
              muxOutConnector[47] = fifoOut[34][7];
              muxOutConnector[48] = fifoOut[35][7];
              muxOutConnector[49] = fifoOut[36][7];
              muxOutConnector[50] = fifoOut[37][7];
              muxOutConnector[51] = fifoOut[38][7];
       end
       17: begin
              muxOutConnector[0] = fifoOut[37][1];
              muxOutConnector[1] = fifoOut[38][1];
              muxOutConnector[2] = fifoOut[39][1];
              muxOutConnector[3] = fifoOut[40][1];
              muxOutConnector[4] = fifoOut[41][1];
              muxOutConnector[5] = fifoOut[42][1];
              muxOutConnector[6] = fifoOut[43][1];
              muxOutConnector[7] = fifoOut[44][1];
              muxOutConnector[8] = fifoOut[45][1];
              muxOutConnector[9] = fifoOut[46][1];
              muxOutConnector[10] = fifoOut[47][1];
              muxOutConnector[11] = fifoOut[48][1];
              muxOutConnector[12] = fifoOut[49][1];
              muxOutConnector[13] = fifoOut[50][1];
              muxOutConnector[14] = fifoOut[51][1];
              muxOutConnector[15] = fifoOut[26][0];
              muxOutConnector[16] = fifoOut[27][0];
              muxOutConnector[17] = fifoOut[28][0];
              muxOutConnector[18] = fifoOut[29][0];
              muxOutConnector[19] = fifoOut[30][0];
              muxOutConnector[20] = fifoOut[31][0];
              muxOutConnector[21] = fifoOut[32][0];
              muxOutConnector[22] = fifoOut[33][0];
              muxOutConnector[23] = fifoOut[34][0];
              muxOutConnector[24] = fifoOut[35][0];
              muxOutConnector[25] = fifoOut[36][0];
              muxOutConnector[26] = fifoOut[39][8];
              muxOutConnector[27] = fifoOut[40][8];
              muxOutConnector[28] = fifoOut[41][8];
              muxOutConnector[29] = fifoOut[42][8];
              muxOutConnector[30] = fifoOut[43][8];
              muxOutConnector[31] = fifoOut[44][8];
              muxOutConnector[32] = fifoOut[45][8];
              muxOutConnector[33] = fifoOut[46][8];
              muxOutConnector[34] = fifoOut[47][8];
              muxOutConnector[35] = fifoOut[48][8];
              muxOutConnector[36] = fifoOut[49][8];
              muxOutConnector[37] = fifoOut[50][8];
              muxOutConnector[38] = fifoOut[51][8];
              muxOutConnector[39] = fifoOut[26][7];
              muxOutConnector[40] = fifoOut[27][7];
              muxOutConnector[41] = fifoOut[28][7];
              muxOutConnector[42] = fifoOut[29][7];
              muxOutConnector[43] = fifoOut[30][7];
              muxOutConnector[44] = fifoOut[31][7];
              muxOutConnector[45] = fifoOut[32][7];
              muxOutConnector[46] = fifoOut[33][7];
              muxOutConnector[47] = fifoOut[34][7];
              muxOutConnector[48] = fifoOut[35][7];
              muxOutConnector[49] = fifoOut[36][7];
              muxOutConnector[50] = fifoOut[37][7];
              muxOutConnector[51] = fifoOut[38][7];
       end
       18: begin
              muxOutConnector[0] = fifoOut[37][1];
              muxOutConnector[1] = fifoOut[38][1];
              muxOutConnector[2] = fifoOut[39][1];
              muxOutConnector[3] = fifoOut[40][1];
              muxOutConnector[4] = fifoOut[41][1];
              muxOutConnector[5] = fifoOut[42][1];
              muxOutConnector[6] = fifoOut[43][1];
              muxOutConnector[7] = fifoOut[44][1];
              muxOutConnector[8] = fifoOut[45][1];
              muxOutConnector[9] = fifoOut[46][1];
              muxOutConnector[10] = fifoOut[47][1];
              muxOutConnector[11] = fifoOut[48][1];
              muxOutConnector[12] = fifoOut[49][1];
              muxOutConnector[13] = fifoOut[50][1];
              muxOutConnector[14] = fifoOut[51][1];
              muxOutConnector[15] = fifoOut[26][0];
              muxOutConnector[16] = fifoOut[27][0];
              muxOutConnector[17] = fifoOut[28][0];
              muxOutConnector[18] = fifoOut[29][0];
              muxOutConnector[19] = fifoOut[30][0];
              muxOutConnector[20] = fifoOut[31][0];
              muxOutConnector[21] = fifoOut[32][0];
              muxOutConnector[22] = fifoOut[33][0];
              muxOutConnector[23] = fifoOut[34][0];
              muxOutConnector[24] = fifoOut[35][0];
              muxOutConnector[25] = fifoOut[36][0];
              muxOutConnector[26] = fifoOut[39][8];
              muxOutConnector[27] = fifoOut[40][8];
              muxOutConnector[28] = fifoOut[41][8];
              muxOutConnector[29] = fifoOut[42][8];
              muxOutConnector[30] = fifoOut[43][8];
              muxOutConnector[31] = fifoOut[44][8];
              muxOutConnector[32] = fifoOut[45][8];
              muxOutConnector[33] = fifoOut[46][8];
              muxOutConnector[34] = fifoOut[47][8];
              muxOutConnector[35] = fifoOut[48][8];
              muxOutConnector[36] = fifoOut[49][8];
              muxOutConnector[37] = fifoOut[50][8];
              muxOutConnector[38] = fifoOut[51][8];
              muxOutConnector[39] = fifoOut[26][7];
              muxOutConnector[40] = fifoOut[27][7];
              muxOutConnector[41] = fifoOut[28][7];
              muxOutConnector[42] = fifoOut[29][7];
              muxOutConnector[43] = fifoOut[30][7];
              muxOutConnector[44] = fifoOut[31][7];
              muxOutConnector[45] = fifoOut[32][7];
              muxOutConnector[46] = fifoOut[33][7];
              muxOutConnector[47] = fifoOut[34][7];
              muxOutConnector[48] = fifoOut[35][7];
              muxOutConnector[49] = fifoOut[36][7];
              muxOutConnector[50] = fifoOut[37][7];
              muxOutConnector[51] = fifoOut[38][7];
       end
       19: begin
              muxOutConnector[0] = fifoOut[37][1];
              muxOutConnector[1] = fifoOut[38][1];
              muxOutConnector[2] = fifoOut[39][1];
              muxOutConnector[3] = fifoOut[40][1];
              muxOutConnector[4] = fifoOut[41][1];
              muxOutConnector[5] = fifoOut[42][1];
              muxOutConnector[6] = fifoOut[43][1];
              muxOutConnector[7] = fifoOut[44][1];
              muxOutConnector[8] = fifoOut[45][1];
              muxOutConnector[9] = fifoOut[46][1];
              muxOutConnector[10] = fifoOut[47][1];
              muxOutConnector[11] = fifoOut[48][1];
              muxOutConnector[12] = fifoOut[49][1];
              muxOutConnector[13] = fifoOut[50][1];
              muxOutConnector[14] = fifoOut[51][1];
              muxOutConnector[15] = fifoOut[26][0];
              muxOutConnector[16] = fifoOut[27][0];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[39][8];
              muxOutConnector[27] = fifoOut[40][8];
              muxOutConnector[28] = fifoOut[41][8];
              muxOutConnector[29] = fifoOut[42][8];
              muxOutConnector[30] = fifoOut[21][7];
              muxOutConnector[31] = fifoOut[22][7];
              muxOutConnector[32] = fifoOut[23][7];
              muxOutConnector[33] = fifoOut[24][7];
              muxOutConnector[34] = fifoOut[25][7];
              muxOutConnector[35] = fifoOut[0][6];
              muxOutConnector[36] = fifoOut[1][6];
              muxOutConnector[37] = fifoOut[2][6];
              muxOutConnector[38] = fifoOut[3][6];
              muxOutConnector[39] = fifoOut[4][6];
              muxOutConnector[40] = fifoOut[5][6];
              muxOutConnector[41] = fifoOut[6][6];
              muxOutConnector[42] = fifoOut[7][6];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
