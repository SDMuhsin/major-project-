`timescale 1ns / 1ps

module ne_funcgenROM(f, romaddress, rden);
parameter Z=511;//circulant size
parameter MB=2;//num of blk columns of G parity part
parameter ADDRESSWIDTH=4;
parameter READDEFAULTCASE = (2**ADDRESSWIDTH)-1;

output reg[(MB*Z)-1:0] f;
input[(ADDRESSWIDTH)-1:0] romaddress;
input rden;

wire[(ADDRESSWIDTH)-1:0] romaddress_case = rden ? romaddress : READDEFAULTCASE;

always@(*)
begin
  case(romaddress_case)
     0: begin
         f=1022'h0AB7EAD98AA507BFDDFD51919FE09C3D7B20CEE21311C4A091ACEA4A84D273C40D1A5B8DF9A5F0457D6D7B2D914EDE926555D378A75A41455390D768C3C86EB39A156B821A62942A8C145DA1E4F708E1512BCFFA61CE44086ABD8E0E9940D0270F3A5C6A02CFB3848D8FBA026807644813C604448FAAE19F4F903A319496174A;
       end
     1: begin
         f=1022'hF62B21CF0AEE0649FA67B7D0EA6551C1CD194CA77501E0FCF8C85867B9CF679C18BCF7939E10F8550661848A4E0A9E9EDB7DAB9EDABA18C168C8E28AACDDEAB18C96E3E90D5AAE24ACC188A2448F6453E002F74C938D822291F6016E101050DE352F20E91A52D4B27F49FA58DAF55EEEA1E18E36635DCB68018FEBAE755E00E2;
       end
     2: begin
         f=1022'hEB40D4728A105EC14A76709F248EB0C041FFDDD4186DAFD7998104C3BEC00FC95AF0388BE2BF3AFB786C39D9F290790F57EBC60B0963114088D1B4EABC87AC94C04DF1DD77F1C20C1FB570D7DD7A1219EAECEA4B2877282651B0FFE713DF338A63263BC0E324A87E2DC1AD64C9F10AAA585ED6905946EE167A73CF04AD2AF921;
       end
     3: begin
         f=1022'h1CD6547FB9BC832408A5B2522000CD179B1549B154648C1153155AE2813F037190B5A0B652D1652D465C0DF7C56D605EC9BC5B428CC0B024E0D04A08BDB4AC8D63B40E7BF93C1C0714789315917A05F9A02DFDC9188D451A684260432323BBA18EDFEEE974151733A15D6B299DA8D95EF701BBF4FB731EE505878EFCBF39EAE6;
       end
     4: begin
         f=1022'h023102AF5C83060E8975C15B4C52BC116F3488103C223ED377CF063A0F7DD7EEC465C0CBEEA5A9E431A736D8B7E415CB71FE2E54FE3ED01CD7EB558788686E6DDD76029801F05D6D703762291091038B0A71A84DAEF383656962A0ED232839D1D3A51DB24B8CF4592FFE50E9873840C77FD106C2C5D4826D260E53D1E51910E4;
       end
     5: begin
         f=1022'h1A60CD1F1C282A1612657E8C7C1420332CA245C0756F78744C807966C3E1326438878BD2CCC83388415A612705AB192B3512EEF0D95248F7B73E5B0F412BF76DEE8696D2F73193E7C90A0591B7B123A14070D32C28DBD7DE23A97066067C0BDB851F011E4BD1E62826BCCCEB6EC116CDEFFE672461048526004BBB8976CB9AF6;
       end
     6: begin
         f=1022'h123B342A892E7EE4026D7C6DF1B307434321011876A7024EF88EC171ABE2A7F12B7500FAB40ECAAA263D0F195BE18547367AE8434F3AA7FEF3577D36BDF478D8BE222975D325A487FE560A6D146311578D9C5501D28BC0A1FB48C9BDA173E869133A3AA9506C42AE9F466E85611FC5F8F74E439638D66D2F00C682987A96D888;
       end
     7: begin
         f=1022'hE3852D7E63A3557F23A6D3B914F1A58F814851EA15EB078219D76668C239C9A7EB158035EC5577A32C6EB1E1BD16D1AD48C1CDA4B79D17F7C41C93768E3F424E800DB8D7FDC08BDE7C5AE80154CFF7524A81E01ACD82B4B1FF29388A073137B7C7E74F94D9B823FCE544F5E73B0202E313BF994832EF90D59DBBCD59F4644AAA;
       end
     8: begin
         f=1022'h034001169D133CBEFCD257B9CD39C7F5B32E3079F5D64F0BA187B395CA2062DA97ACB4540D974FE9C98950107359502024686C91DD51B77448C94D1C22B567E82BD6DFF9A022843A90BFBC3B66D06483E0808C217041BEEF07D5AD59E85095C086F17F69832E816C23EB5B70EC1040A562131F33783958D1F592779B773BAC32;
       end
     9: begin
         f=1022'hF595E9B2B33EF82D0E64AA2226D6A0ADCD179D5932EE1CF401B336449D0FF775754CA56650716E61A43F963D59865C7F017F53830514306649822CAA72C152F698459B02819146FBC1A04C24B3EC7545484151F03FD96CC3B74B8C5BED902F694C3A5783E0D14A1BFA1D51FC37A70EC020C5C44ED4930F4334E168C18A9E42BC;
       end
    10: begin
         f=1022'hFF08378FF9248C979757831A447133F774CA73BB04CAE27D37FD072120C12D3FADB2E3A7D8B5626448DE004699D6A7FCBA91F72DE8A09348B702817F97C7250397865287840D00243278F41CE1156D1868F24E02F91D3A1886ACE906CE741662B40B4EFDFB90F76C1ADD884D920AFA8B3427EEB84A759FA02E00635743F50B94;
       end
    11: begin
         f=1022'hFB71042768A893906C7CDD59148A660752DFA230DA84B6AD93A471D93310F33B0623B231615723FD222EE4400D80AFBD0F6FB12988412241A8B37176F5040D0C2F910C2F1DE383B5D28D56B58CCE46305E6B874122DC3A49389B736C6EA93EF8349EE0850E4728DADF49FFBA9C7D09C599AB9C7A18A9B0D5FC639DFA02C9D711;
       end
    12: begin
         f=1022'hF97245108AEEB44C4A0B68E511C0CB647694DAF15F7BB646AD67258D25DEAD46B569544EECFBCE5E0B18C9088AF92B5199BA1DE44B574AD6ECAF6FE1D28FB82FCD2498C31BDE61E39433D6AF4D4E9BB602FAB31C5A45E7A95D0D7911046F1F55984DB7EA60C067CD10F7A393182502F138C773AB54535D56BE5698896175A55C;
       end
    13: begin
         f=1022'h1BDB7273E8342918E097B1C1F5FEF32A150AEF5E11184782B5BD5A1D8071E94578B0AC722D7BF49E8C78D391294371FFBA7B88FABF8CC03A62B940CE60D669DFD73E10FD424084F2660E08B6507AE60BD27B1EE8E4A069CEFA4BA7FE0875B8BF16B630DB6E152D1502D06BDF6AEB2A5D5CFD49CEDBE1ABE12EB21C34552F004A;
       end
    default: begin
               f=0;
             end
  endcase
end
endmodule
