`timescale 1ns / 1ps

module ne_testcodestimulusROM(dout, rd_address, rd_en);
parameter DEPTH=257;//(8160+64)/32
parameter ADDRESSWIDTH=9;//ceil(log2(DEPTH))
parameter W=6;
parameter DW=192;//32xW
parameter READDEFAULTCASE=9'b1_1111_1111;

output reg[DW-1:0] dout;
input[ADDRESSWIDTH-1:0] rd_address;
input rd_en;

wire[ADDRESSWIDTH-1:0] rd_address_case;
assign rd_address_case = rd_en ? rd_address : READDEFAULTCASE;
always@(*) begin
 case(rd_address_case)
   0: begin
        dout = {6'b110111, 6'b000111, 6'b001011, 6'b001011, 6'b110110, 6'b110101, 6'b111000, 6'b001010, 6'b000000, 6'b110010, 6'b111101, 6'b110011, 6'b111010, 6'b001110, 6'b110111, 6'b110100, 6'b111111, 6'b111000, 6'b111011, 6'b001001, 6'b110111, 6'b111010, 6'b001010, 6'b111100, 6'b111010, 6'b110111, 6'b111010, 6'b001001, 6'b000110, 6'b000100, 6'b111101, 6'b000011};
      end
   1: begin
        dout = {6'b001110, 6'b000111, 6'b000101, 6'b001001, 6'b001111, 6'b111001, 6'b111110, 6'b110100, 6'b111101, 6'b111010, 6'b110111, 6'b111010, 6'b110110, 6'b001000, 6'b010011, 6'b000001, 6'b000001, 6'b110100, 6'b001001, 6'b001100, 6'b110110, 6'b000001, 6'b001011, 6'b001101, 6'b001001, 6'b110100, 6'b001010, 6'b001001, 6'b110110, 6'b001101, 6'b001000, 6'b111001};
      end
   2: begin
        dout = {6'b111010, 6'b001011, 6'b110100, 6'b001111, 6'b110101, 6'b110110, 6'b001010, 6'b001110, 6'b001011, 6'b111101, 6'b001000, 6'b111011, 6'b001110, 6'b000100, 6'b001001, 6'b101110, 6'b111010, 6'b001010, 6'b000010, 6'b110111, 6'b000100, 6'b111000, 6'b110101, 6'b000110, 6'b000101, 6'b110110, 6'b001110, 6'b000111, 6'b111001, 6'b111101, 6'b001100, 6'b001000};
      end
   3: begin
        dout = {6'b110111, 6'b111001, 6'b110111, 6'b110111, 6'b111000, 6'b111001, 6'b110111, 6'b000011, 6'b110001, 6'b111010, 6'b001101, 6'b111010, 6'b001001, 6'b001000, 6'b111000, 6'b110110, 6'b111000, 6'b110100, 6'b110000, 6'b101111, 6'b110101, 6'b001011, 6'b001000, 6'b110110, 6'b000101, 6'b001001, 6'b001011, 6'b000111, 6'b001011, 6'b111000, 6'b001100, 6'b111001};
      end
   4: begin
        dout = {6'b000100, 6'b000100, 6'b001100, 6'b111001, 6'b110111, 6'b111011, 6'b010001, 6'b110111, 6'b111000, 6'b000101, 6'b110110, 6'b000101, 6'b001001, 6'b000010, 6'b110101, 6'b001100, 6'b001010, 6'b111001, 6'b000111, 6'b111000, 6'b110111, 6'b001001, 6'b110010, 6'b111100, 6'b000111, 6'b111001, 6'b001001, 6'b110111, 6'b111101, 6'b001000, 6'b111001, 6'b000111};
      end
   5: begin
        dout = {6'b010000, 6'b000010, 6'b111011, 6'b110011, 6'b110110, 6'b111110, 6'b110111, 6'b001000, 6'b000011, 6'b110111, 6'b111111, 6'b111001, 6'b110101, 6'b110101, 6'b001100, 6'b110110, 6'b110101, 6'b001001, 6'b001110, 6'b000100, 6'b110100, 6'b001000, 6'b110110, 6'b001000, 6'b001111, 6'b110001, 6'b110000, 6'b000100, 6'b110101, 6'b010000, 6'b000010, 6'b000001};
      end
   6: begin
        dout = {6'b110110, 6'b110111, 6'b111110, 6'b111010, 6'b111001, 6'b111100, 6'b110100, 6'b001100, 6'b000000, 6'b110110, 6'b001010, 6'b111000, 6'b001010, 6'b111010, 6'b000000, 6'b110011, 6'b110111, 6'b111000, 6'b111010, 6'b000001, 6'b001101, 6'b111010, 6'b001100, 6'b000001, 6'b000110, 6'b110101, 6'b110100, 6'b110110, 6'b111100, 6'b001011, 6'b000101, 6'b111010};
      end
   7: begin
        dout = {6'b001110, 6'b001000, 6'b111010, 6'b000111, 6'b110101, 6'b110011, 6'b001010, 6'b111010, 6'b001000, 6'b110101, 6'b000110, 6'b000000, 6'b111001, 6'b110110, 6'b000111, 6'b000101, 6'b110010, 6'b000110, 6'b000100, 6'b111110, 6'b001011, 6'b110111, 6'b000100, 6'b110010, 6'b110110, 6'b110010, 6'b001100, 6'b110100, 6'b000001, 6'b000100, 6'b110011, 6'b000100};
      end
   8: begin
        dout = {6'b111001, 6'b000010, 6'b110111, 6'b110101, 6'b000001, 6'b111010, 6'b111000, 6'b001100, 6'b111010, 6'b110111, 6'b110110, 6'b001001, 6'b111110, 6'b110111, 6'b000101, 6'b110111, 6'b110111, 6'b001010, 6'b110110, 6'b010001, 6'b000001, 6'b111000, 6'b110011, 6'b111001, 6'b111111, 6'b000110, 6'b111111, 6'b111001, 6'b110000, 6'b110110, 6'b111101, 6'b111101};
      end
   9: begin
        dout = {6'b110111, 6'b111010, 6'b000111, 6'b110101, 6'b001111, 6'b110101, 6'b000101, 6'b000000, 6'b000110, 6'b111000, 6'b000011, 6'b110110, 6'b110111, 6'b001010, 6'b111110, 6'b000011, 6'b111001, 6'b000010, 6'b111010, 6'b001011, 6'b001010, 6'b001010, 6'b111100, 6'b001000, 6'b111010, 6'b000110, 6'b110010, 6'b000010, 6'b001010, 6'b110011, 6'b001110, 6'b110101};
      end
   10: begin
        dout = {6'b001010, 6'b000011, 6'b000010, 6'b001100, 6'b111010, 6'b110011, 6'b001000, 6'b111010, 6'b110011, 6'b000100, 6'b110111, 6'b001011, 6'b110010, 6'b110111, 6'b000010, 6'b110111, 6'b111001, 6'b110011, 6'b110111, 6'b001010, 6'b001011, 6'b000110, 6'b111011, 6'b111011, 6'b111111, 6'b111000, 6'b110011, 6'b000101, 6'b001000, 6'b110101, 6'b110111, 6'b111001};
      end
   11: begin
        dout = {6'b110110, 6'b001010, 6'b001010, 6'b110010, 6'b101111, 6'b111000, 6'b110100, 6'b001001, 6'b110100, 6'b000101, 6'b001000, 6'b111000, 6'b111000, 6'b000011, 6'b111100, 6'b111110, 6'b001010, 6'b001010, 6'b111001, 6'b110111, 6'b111100, 6'b110111, 6'b110110, 6'b000100, 6'b110110, 6'b111011, 6'b111000, 6'b000011, 6'b001010, 6'b111110, 6'b110110, 6'b111101};
      end
   12: begin
        dout = {6'b000101, 6'b110101, 6'b001011, 6'b000101, 6'b000010, 6'b000010, 6'b111100, 6'b110111, 6'b111011, 6'b111011, 6'b001010, 6'b001001, 6'b110101, 6'b010001, 6'b001000, 6'b110111, 6'b110100, 6'b110110, 6'b111101, 6'b000000, 6'b110101, 6'b000100, 6'b110100, 6'b111010, 6'b001010, 6'b110101, 6'b000101, 6'b000110, 6'b000000, 6'b000111, 6'b110011, 6'b000101};
      end
   13: begin
        dout = {6'b000011, 6'b000011, 6'b000100, 6'b111011, 6'b110110, 6'b001001, 6'b111000, 6'b001101, 6'b000100, 6'b110111, 6'b000001, 6'b000111, 6'b000110, 6'b111010, 6'b000010, 6'b000101, 6'b111111, 6'b110100, 6'b110111, 6'b110101, 6'b000110, 6'b111100, 6'b000010, 6'b001011, 6'b111100, 6'b111000, 6'b000010, 6'b000111, 6'b000001, 6'b000100, 6'b111100, 6'b111000};
      end
   14: begin
        dout = {6'b111001, 6'b001001, 6'b111010, 6'b111000, 6'b110011, 6'b001001, 6'b110010, 6'b001000, 6'b111001, 6'b000100, 6'b000110, 6'b001100, 6'b110100, 6'b110100, 6'b001000, 6'b111111, 6'b111110, 6'b110110, 6'b110111, 6'b111110, 6'b110011, 6'b000011, 6'b001001, 6'b000110, 6'b001110, 6'b111010, 6'b000111, 6'b110111, 6'b111101, 6'b000110, 6'b110100, 6'b110101};
      end
   15: begin
        dout = {6'b010000, 6'b000111, 6'b110100, 6'b110011, 6'b001000, 6'b001011, 6'b001100, 6'b110110, 6'b110001, 6'b111010, 6'b000101, 6'b000111, 6'b111000, 6'b110110, 6'b001001, 6'b111000, 6'b000100, 6'b110010, 6'b110100, 6'b001001, 6'b110010, 6'b000010, 6'b110010, 6'b110011, 6'b000110, 6'b001000, 6'b110111, 6'b000101, 6'b111000, 6'b001010, 6'b001000, 6'b110111};
      end
   16: begin
        dout = {6'b111100, 6'b000110, 6'b000011, 6'b110111, 6'b001010, 6'b001100, 6'b111011, 6'b000011, 6'b001100, 6'b110110, 6'b110101, 6'b000000, 6'b000111, 6'b001011, 6'b111101, 6'b111100, 6'b111001, 6'b000111, 6'b000110, 6'b110101, 6'b111011, 6'b001010, 6'b110010, 6'b110011, 6'b110101, 6'b000111, 6'b000111, 6'b001010, 6'b000011, 6'b110011, 6'b110110, 6'b110011};
      end
   17: begin
        dout = {6'b110110, 6'b101111, 6'b000100, 6'b111011, 6'b111001, 6'b001001, 6'b110011, 6'b110111, 6'b110011, 6'b110111, 6'b001010, 6'b001100, 6'b000111, 6'b111101, 6'b110000, 6'b110111, 6'b111001, 6'b001010, 6'b001010, 6'b111001, 6'b000111, 6'b001000, 6'b110101, 6'b110010, 6'b010000, 6'b111010, 6'b000010, 6'b110101, 6'b000100, 6'b000111, 6'b110100, 6'b111100};
      end
   18: begin
        dout = {6'b110101, 6'b000011, 6'b000101, 6'b001000, 6'b110110, 6'b001001, 6'b001101, 6'b111001, 6'b000111, 6'b110010, 6'b111101, 6'b001001, 6'b001010, 6'b000101, 6'b111000, 6'b001011, 6'b111111, 6'b110111, 6'b001101, 6'b110011, 6'b001000, 6'b000110, 6'b110111, 6'b001111, 6'b111010, 6'b101111, 6'b111100, 6'b110010, 6'b111000, 6'b110101, 6'b001001, 6'b111000};
      end
   19: begin
        dout = {6'b111100, 6'b000001, 6'b000111, 6'b000101, 6'b110110, 6'b111101, 6'b110100, 6'b001101, 6'b010001, 6'b110110, 6'b111011, 6'b111111, 6'b001000, 6'b110111, 6'b000110, 6'b110010, 6'b010000, 6'b001011, 6'b000101, 6'b111001, 6'b000110, 6'b111000, 6'b111110, 6'b001111, 6'b001001, 6'b001100, 6'b001001, 6'b110110, 6'b110111, 6'b110001, 6'b110100, 6'b000010};
      end
   20: begin
        dout = {6'b000101, 6'b000101, 6'b000011, 6'b110100, 6'b110100, 6'b110110, 6'b001101, 6'b111001, 6'b000111, 6'b111001, 6'b000011, 6'b111100, 6'b000010, 6'b000110, 6'b000111, 6'b110100, 6'b111011, 6'b001011, 6'b001110, 6'b001010, 6'b001010, 6'b111110, 6'b110111, 6'b001000, 6'b001100, 6'b000110, 6'b111000, 6'b000000, 6'b001001, 6'b111000, 6'b110111, 6'b110001};
      end
   21: begin
        dout = {6'b001011, 6'b110100, 6'b000110, 6'b000111, 6'b001010, 6'b001100, 6'b111001, 6'b001001, 6'b111010, 6'b000111, 6'b001100, 6'b110001, 6'b111100, 6'b110110, 6'b111000, 6'b110111, 6'b110110, 6'b110011, 6'b111010, 6'b111001, 6'b110101, 6'b000111, 6'b111010, 6'b110010, 6'b001000, 6'b000000, 6'b001101, 6'b000000, 6'b001010, 6'b001010, 6'b110010, 6'b001101};
      end
   22: begin
        dout = {6'b111010, 6'b001001, 6'b001000, 6'b111011, 6'b110011, 6'b001001, 6'b000111, 6'b001001, 6'b001100, 6'b000011, 6'b111000, 6'b110101, 6'b111110, 6'b110101, 6'b000100, 6'b110111, 6'b101110, 6'b110100, 6'b111100, 6'b111010, 6'b000010, 6'b000110, 6'b110110, 6'b000101, 6'b000110, 6'b111000, 6'b000110, 6'b000101, 6'b000000, 6'b110010, 6'b001010, 6'b101111};
      end
   23: begin
        dout = {6'b110000, 6'b110010, 6'b111001, 6'b110100, 6'b101111, 6'b000011, 6'b001111, 6'b111000, 6'b000010, 6'b110001, 6'b000111, 6'b111110, 6'b001011, 6'b110101, 6'b001011, 6'b000110, 6'b001100, 6'b111011, 6'b110000, 6'b110101, 6'b000100, 6'b001000, 6'b111011, 6'b110111, 6'b111000, 6'b001000, 6'b001000, 6'b001011, 6'b111101, 6'b111101, 6'b001011, 6'b000011};
      end
   24: begin
        dout = {6'b111001, 6'b000110, 6'b001010, 6'b110100, 6'b001000, 6'b001001, 6'b110001, 6'b111001, 6'b110011, 6'b000101, 6'b110101, 6'b110101, 6'b000000, 6'b111101, 6'b001100, 6'b000101, 6'b001011, 6'b111001, 6'b110111, 6'b110011, 6'b111100, 6'b000000, 6'b000110, 6'b110101, 6'b110010, 6'b111010, 6'b111001, 6'b000101, 6'b001010, 6'b001101, 6'b000100, 6'b000111};
      end
   25: begin
        dout = {6'b110110, 6'b000110, 6'b111000, 6'b111000, 6'b111001, 6'b110001, 6'b111000, 6'b110110, 6'b001001, 6'b000101, 6'b110100, 6'b001101, 6'b111010, 6'b001000, 6'b001011, 6'b000101, 6'b111010, 6'b110111, 6'b111000, 6'b001100, 6'b110101, 6'b111111, 6'b001011, 6'b110111, 6'b111101, 6'b001011, 6'b001000, 6'b111010, 6'b001000, 6'b110111, 6'b111010, 6'b000001};
      end
   26: begin
        dout = {6'b110010, 6'b000010, 6'b001111, 6'b111000, 6'b001000, 6'b111011, 6'b001100, 6'b111000, 6'b001011, 6'b001101, 6'b111010, 6'b000000, 6'b000101, 6'b000101, 6'b111101, 6'b110111, 6'b110101, 6'b110101, 6'b001100, 6'b001110, 6'b111000, 6'b001010, 6'b110111, 6'b000110, 6'b001000, 6'b001101, 6'b000011, 6'b111011, 6'b111001, 6'b000101, 6'b110011, 6'b110011};
      end
   27: begin
        dout = {6'b000100, 6'b110010, 6'b110101, 6'b001000, 6'b000101, 6'b001100, 6'b001011, 6'b110100, 6'b010011, 6'b001000, 6'b110101, 6'b110101, 6'b000110, 6'b001001, 6'b001001, 6'b111011, 6'b001000, 6'b111001, 6'b111010, 6'b000010, 6'b001000, 6'b001110, 6'b000111, 6'b110001, 6'b001010, 6'b000100, 6'b110011, 6'b001001, 6'b111011, 6'b001000, 6'b111000, 6'b110110};
      end
   28: begin
        dout = {6'b110111, 6'b000101, 6'b111000, 6'b110111, 6'b000011, 6'b001110, 6'b111100, 6'b110101, 6'b000110, 6'b000111, 6'b000111, 6'b001101, 6'b000111, 6'b001000, 6'b000111, 6'b110010, 6'b110100, 6'b000010, 6'b000100, 6'b000111, 6'b110011, 6'b110100, 6'b111110, 6'b000110, 6'b111100, 6'b010000, 6'b000110, 6'b001111, 6'b111101, 6'b110111, 6'b110111, 6'b110100};
      end
   29: begin
        dout = {6'b111000, 6'b111001, 6'b001011, 6'b001000, 6'b000101, 6'b000111, 6'b111100, 6'b000101, 6'b110000, 6'b110011, 6'b000110, 6'b001100, 6'b111010, 6'b001100, 6'b000101, 6'b001010, 6'b110010, 6'b101100, 6'b001111, 6'b110111, 6'b001011, 6'b110111, 6'b001100, 6'b000110, 6'b001000, 6'b000101, 6'b111000, 6'b111101, 6'b110111, 6'b111100, 6'b000100, 6'b000100};
      end
   30: begin
        dout = {6'b001101, 6'b110100, 6'b110110, 6'b001001, 6'b110101, 6'b110011, 6'b000100, 6'b111010, 6'b001011, 6'b001001, 6'b110111, 6'b111011, 6'b000111, 6'b110001, 6'b000101, 6'b111001, 6'b001100, 6'b110011, 6'b111011, 6'b001001, 6'b000111, 6'b111000, 6'b111010, 6'b001011, 6'b001000, 6'b111011, 6'b111010, 6'b000110, 6'b001010, 6'b110110, 6'b111011, 6'b111010};
      end
   31: begin
        dout = {6'b111011, 6'b110010, 6'b111010, 6'b111100, 6'b000000, 6'b001101, 6'b110010, 6'b110111, 6'b000110, 6'b111001, 6'b000110, 6'b110101, 6'b000000, 6'b110110, 6'b000010, 6'b110110, 6'b000100, 6'b110110, 6'b111010, 6'b111001, 6'b111001, 6'b111010, 6'b000111, 6'b001011, 6'b110110, 6'b111011, 6'b110010, 6'b110011, 6'b000101, 6'b001000, 6'b001100, 6'b000111};
      end
   32: begin
        dout = {6'b111101, 6'b000001, 6'b110011, 6'b001010, 6'b000101, 6'b001010, 6'b110101, 6'b000001, 6'b001001, 6'b000111, 6'b111010, 6'b110100, 6'b110010, 6'b111011, 6'b001001, 6'b000111, 6'b111111, 6'b000100, 6'b110111, 6'b001011, 6'b000011, 6'b001011, 6'b001011, 6'b001000, 6'b111011, 6'b111101, 6'b111010, 6'b110111, 6'b111010, 6'b000110, 6'b001110, 6'b001010};
      end
   33: begin
        dout = {6'b001110, 6'b001011, 6'b111010, 6'b110111, 6'b110111, 6'b000110, 6'b110111, 6'b111010, 6'b111000, 6'b111111, 6'b111000, 6'b110101, 6'b111000, 6'b110110, 6'b001011, 6'b000101, 6'b000110, 6'b111000, 6'b111100, 6'b110010, 6'b000101, 6'b110001, 6'b000000, 6'b001000, 6'b110111, 6'b000101, 6'b101111, 6'b110111, 6'b000010, 6'b111000, 6'b110110, 6'b000001};
      end
   34: begin
        dout = {6'b111111, 6'b001001, 6'b111100, 6'b110010, 6'b001101, 6'b110010, 6'b000110, 6'b110110, 6'b111010, 6'b110110, 6'b000101, 6'b000011, 6'b001010, 6'b110100, 6'b110010, 6'b110101, 6'b001101, 6'b110100, 6'b001001, 6'b000101, 6'b001010, 6'b001111, 6'b001000, 6'b000011, 6'b110000, 6'b111010, 6'b000001, 6'b000011, 6'b111001, 6'b110110, 6'b111000, 6'b111000};
      end
   35: begin
        dout = {6'b000110, 6'b000111, 6'b000101, 6'b111000, 6'b000010, 6'b001101, 6'b001000, 6'b001110, 6'b001001, 6'b111011, 6'b111010, 6'b110100, 6'b111000, 6'b000101, 6'b110001, 6'b111101, 6'b110101, 6'b000000, 6'b110011, 6'b000101, 6'b001010, 6'b001100, 6'b111000, 6'b111010, 6'b110111, 6'b000011, 6'b000011, 6'b111100, 6'b110111, 6'b001000, 6'b001110, 6'b000011};
      end
   36: begin
        dout = {6'b110111, 6'b110010, 6'b110111, 6'b111001, 6'b110011, 6'b001110, 6'b110100, 6'b000000, 6'b000110, 6'b001000, 6'b110101, 6'b001000, 6'b111010, 6'b000110, 6'b001100, 6'b110110, 6'b110101, 6'b001100, 6'b101110, 6'b110001, 6'b111011, 6'b000100, 6'b001010, 6'b111001, 6'b111100, 6'b111001, 6'b001001, 6'b001011, 6'b010011, 6'b111001, 6'b111010, 6'b110011};
      end
   37: begin
        dout = {6'b110111, 6'b111001, 6'b000111, 6'b111000, 6'b111001, 6'b110100, 6'b110101, 6'b000110, 6'b111011, 6'b000110, 6'b001000, 6'b000111, 6'b001100, 6'b001100, 6'b111001, 6'b000101, 6'b001110, 6'b001000, 6'b110011, 6'b000111, 6'b111001, 6'b111010, 6'b000000, 6'b000110, 6'b001000, 6'b110100, 6'b111010, 6'b111011, 6'b110110, 6'b000001, 6'b000110, 6'b001101};
      end
   38: begin
        dout = {6'b111001, 6'b111010, 6'b000110, 6'b110100, 6'b000111, 6'b001001, 6'b111010, 6'b111000, 6'b001000, 6'b001001, 6'b000110, 6'b000111, 6'b000001, 6'b000111, 6'b000111, 6'b110001, 6'b111010, 6'b111001, 6'b110101, 6'b000011, 6'b000100, 6'b001100, 6'b010001, 6'b000110, 6'b001010, 6'b110110, 6'b111001, 6'b111000, 6'b110111, 6'b110110, 6'b111001, 6'b001100};
      end
   39: begin
        dout = {6'b111011, 6'b111111, 6'b001101, 6'b001011, 6'b001001, 6'b111100, 6'b110100, 6'b111011, 6'b111010, 6'b111001, 6'b111001, 6'b111011, 6'b000100, 6'b111110, 6'b000100, 6'b000110, 6'b111010, 6'b001000, 6'b110000, 6'b111001, 6'b000110, 6'b110101, 6'b001001, 6'b110101, 6'b110110, 6'b000100, 6'b001001, 6'b110011, 6'b000111, 6'b110001, 6'b001011, 6'b001010};
      end
   40: begin
        dout = {6'b001010, 6'b110111, 6'b111000, 6'b000101, 6'b111000, 6'b111001, 6'b110011, 6'b110110, 6'b000101, 6'b111011, 6'b111000, 6'b111000, 6'b000011, 6'b111011, 6'b111010, 6'b110100, 6'b110101, 6'b000101, 6'b000101, 6'b111000, 6'b110111, 6'b000001, 6'b111101, 6'b000101, 6'b111100, 6'b000110, 6'b001001, 6'b111010, 6'b000110, 6'b110110, 6'b111100, 6'b110111};
      end
   41: begin
        dout = {6'b001101, 6'b110011, 6'b110110, 6'b001000, 6'b001000, 6'b001010, 6'b000011, 6'b110110, 6'b111011, 6'b000011, 6'b000010, 6'b000110, 6'b000101, 6'b000111, 6'b000101, 6'b110111, 6'b000110, 6'b000101, 6'b000100, 6'b000101, 6'b111010, 6'b000111, 6'b001001, 6'b001001, 6'b111011, 6'b001110, 6'b111100, 6'b111111, 6'b001001, 6'b000011, 6'b000111, 6'b110111};
      end
   42: begin
        dout = {6'b001000, 6'b111000, 6'b010010, 6'b001001, 6'b001001, 6'b001001, 6'b001100, 6'b000110, 6'b000100, 6'b001011, 6'b111101, 6'b000111, 6'b111011, 6'b000010, 6'b110100, 6'b110111, 6'b110111, 6'b110010, 6'b000010, 6'b111110, 6'b111010, 6'b110110, 6'b000001, 6'b000110, 6'b000111, 6'b110100, 6'b110110, 6'b000111, 6'b110100, 6'b111001, 6'b000101, 6'b001000};
      end
   43: begin
        dout = {6'b111010, 6'b000110, 6'b111010, 6'b111101, 6'b000110, 6'b110111, 6'b110111, 6'b001101, 6'b111011, 6'b001000, 6'b000100, 6'b001000, 6'b111100, 6'b000111, 6'b000111, 6'b001010, 6'b001100, 6'b001010, 6'b001000, 6'b111010, 6'b110001, 6'b001100, 6'b001000, 6'b000100, 6'b001001, 6'b111000, 6'b000111, 6'b110100, 6'b001011, 6'b000100, 6'b111111, 6'b001111};
      end
   44: begin
        dout = {6'b111000, 6'b111010, 6'b001001, 6'b000001, 6'b110111, 6'b000100, 6'b110001, 6'b111110, 6'b000111, 6'b110111, 6'b111010, 6'b000100, 6'b000100, 6'b111001, 6'b110100, 6'b000111, 6'b001010, 6'b111001, 6'b000011, 6'b001010, 6'b001010, 6'b111110, 6'b000110, 6'b111001, 6'b110001, 6'b110110, 6'b111100, 6'b111001, 6'b110001, 6'b001010, 6'b000100, 6'b111000};
      end
   45: begin
        dout = {6'b001000, 6'b001010, 6'b001001, 6'b110011, 6'b001011, 6'b000001, 6'b000110, 6'b001010, 6'b001001, 6'b001010, 6'b111011, 6'b000110, 6'b111011, 6'b110111, 6'b110111, 6'b000100, 6'b111101, 6'b110000, 6'b110111, 6'b111001, 6'b110111, 6'b001001, 6'b001101, 6'b111001, 6'b000110, 6'b111001, 6'b010000, 6'b001010, 6'b000100, 6'b110110, 6'b000111, 6'b001001};
      end
   46: begin
        dout = {6'b110100, 6'b001001, 6'b001001, 6'b111001, 6'b111011, 6'b111011, 6'b111100, 6'b001000, 6'b000010, 6'b110101, 6'b110000, 6'b001110, 6'b111010, 6'b001110, 6'b000110, 6'b111100, 6'b000001, 6'b001001, 6'b001000, 6'b001001, 6'b001010, 6'b110001, 6'b001010, 6'b111110, 6'b111000, 6'b001000, 6'b111001, 6'b111011, 6'b111100, 6'b110111, 6'b000111, 6'b000111};
      end
   47: begin
        dout = {6'b111011, 6'b001001, 6'b111100, 6'b000010, 6'b110100, 6'b111010, 6'b000111, 6'b000110, 6'b001001, 6'b111001, 6'b001101, 6'b110101, 6'b111011, 6'b111111, 6'b111011, 6'b110101, 6'b001011, 6'b001100, 6'b001010, 6'b110110, 6'b110111, 6'b110011, 6'b111101, 6'b110111, 6'b110110, 6'b111010, 6'b110111, 6'b111111, 6'b000100, 6'b111000, 6'b001010, 6'b000111};
      end
   48: begin
        dout = {6'b110000, 6'b001110, 6'b110110, 6'b111000, 6'b000101, 6'b110101, 6'b001100, 6'b001011, 6'b001001, 6'b111001, 6'b110001, 6'b001001, 6'b000100, 6'b110100, 6'b001001, 6'b110111, 6'b001101, 6'b111000, 6'b110110, 6'b001001, 6'b000101, 6'b110010, 6'b111100, 6'b111100, 6'b111000, 6'b000011, 6'b111011, 6'b101110, 6'b000100, 6'b000111, 6'b110001, 6'b110100};
      end
   49: begin
        dout = {6'b110010, 6'b001100, 6'b000101, 6'b000111, 6'b111001, 6'b000101, 6'b111101, 6'b000110, 6'b111000, 6'b001000, 6'b110111, 6'b111110, 6'b110001, 6'b111110, 6'b111010, 6'b000111, 6'b111001, 6'b000110, 6'b110010, 6'b000101, 6'b110110, 6'b001010, 6'b000011, 6'b110010, 6'b001001, 6'b111001, 6'b111011, 6'b111001, 6'b111111, 6'b000110, 6'b111100, 6'b001110};
      end
   50: begin
        dout = {6'b001010, 6'b000111, 6'b000100, 6'b110011, 6'b111100, 6'b111001, 6'b001001, 6'b110110, 6'b111010, 6'b111000, 6'b110100, 6'b001000, 6'b001000, 6'b110010, 6'b111100, 6'b111010, 6'b001000, 6'b110110, 6'b001111, 6'b000111, 6'b000000, 6'b001000, 6'b111001, 6'b111000, 6'b111100, 6'b110100, 6'b110100, 6'b110110, 6'b001110, 6'b001001, 6'b001111, 6'b111010};
      end
   51: begin
        dout = {6'b110000, 6'b110111, 6'b111010, 6'b000110, 6'b111001, 6'b110100, 6'b111010, 6'b110000, 6'b111000, 6'b111011, 6'b110101, 6'b111010, 6'b111010, 6'b110101, 6'b110101, 6'b000100, 6'b000100, 6'b001001, 6'b010001, 6'b111000, 6'b111000, 6'b110011, 6'b110100, 6'b111000, 6'b111110, 6'b000100, 6'b000011, 6'b001000, 6'b110111, 6'b001001, 6'b111101, 6'b000110};
      end
   52: begin
        dout = {6'b111001, 6'b111001, 6'b001000, 6'b111001, 6'b001110, 6'b001001, 6'b000111, 6'b110110, 6'b001000, 6'b111011, 6'b001100, 6'b110010, 6'b110101, 6'b010011, 6'b001100, 6'b111010, 6'b110001, 6'b111000, 6'b000100, 6'b110111, 6'b110011, 6'b111000, 6'b001110, 6'b000011, 6'b001001, 6'b111100, 6'b111000, 6'b001101, 6'b111110, 6'b000101, 6'b001111, 6'b001001};
      end
   53: begin
        dout = {6'b110111, 6'b111100, 6'b110011, 6'b000001, 6'b000101, 6'b110110, 6'b000101, 6'b000110, 6'b110101, 6'b111111, 6'b110111, 6'b111000, 6'b001001, 6'b110011, 6'b000100, 6'b000001, 6'b000101, 6'b000110, 6'b110101, 6'b001011, 6'b000101, 6'b001000, 6'b111001, 6'b000010, 6'b110111, 6'b110010, 6'b110101, 6'b110110, 6'b110101, 6'b110011, 6'b111011, 6'b111001};
      end
   54: begin
        dout = {6'b000110, 6'b000110, 6'b111101, 6'b111100, 6'b110001, 6'b001001, 6'b110011, 6'b001010, 6'b110111, 6'b000111, 6'b111001, 6'b111000, 6'b000111, 6'b111000, 6'b000101, 6'b111001, 6'b111001, 6'b001000, 6'b110100, 6'b001011, 6'b111011, 6'b110100, 6'b111000, 6'b000010, 6'b000000, 6'b110100, 6'b001001, 6'b000101, 6'b111011, 6'b110111, 6'b001010, 6'b111001};
      end
   55: begin
        dout = {6'b110110, 6'b000011, 6'b110111, 6'b111010, 6'b001101, 6'b110111, 6'b001011, 6'b000001, 6'b111001, 6'b111001, 6'b110111, 6'b000101, 6'b000110, 6'b001001, 6'b111101, 6'b110101, 6'b110100, 6'b111101, 6'b110111, 6'b110101, 6'b110001, 6'b000110, 6'b111001, 6'b111010, 6'b000000, 6'b001000, 6'b111001, 6'b110101, 6'b001000, 6'b110110, 6'b000111, 6'b110110};
      end
   56: begin
        dout = {6'b111000, 6'b000101, 6'b110110, 6'b001100, 6'b110100, 6'b000100, 6'b111000, 6'b000011, 6'b111010, 6'b111010, 6'b111000, 6'b000111, 6'b001001, 6'b001000, 6'b001010, 6'b001101, 6'b111001, 6'b000010, 6'b111100, 6'b000110, 6'b111000, 6'b110100, 6'b001001, 6'b000001, 6'b110110, 6'b001011, 6'b110101, 6'b001001, 6'b001001, 6'b000101, 6'b110111, 6'b000111};
      end
   57: begin
        dout = {6'b110101, 6'b101110, 6'b110111, 6'b111011, 6'b001000, 6'b110010, 6'b111100, 6'b000111, 6'b111001, 6'b111011, 6'b000100, 6'b110110, 6'b001001, 6'b000100, 6'b001011, 6'b001001, 6'b001010, 6'b000110, 6'b111001, 6'b001101, 6'b001011, 6'b000011, 6'b110100, 6'b111010, 6'b110100, 6'b000100, 6'b110110, 6'b001001, 6'b111010, 6'b000111, 6'b111001, 6'b001001};
      end
   58: begin
        dout = {6'b111100, 6'b111001, 6'b110111, 6'b110101, 6'b000111, 6'b111010, 6'b110111, 6'b110111, 6'b111010, 6'b000111, 6'b000110, 6'b110001, 6'b000011, 6'b110110, 6'b000101, 6'b110101, 6'b110111, 6'b111000, 6'b111011, 6'b000111, 6'b110100, 6'b111110, 6'b110100, 6'b001000, 6'b000110, 6'b110100, 6'b001101, 6'b001010, 6'b111100, 6'b000011, 6'b110110, 6'b111100};
      end
   59: begin
        dout = {6'b111001, 6'b111000, 6'b001010, 6'b110101, 6'b001000, 6'b001010, 6'b111000, 6'b111001, 6'b001101, 6'b110101, 6'b000000, 6'b110110, 6'b110101, 6'b000110, 6'b000101, 6'b000110, 6'b111101, 6'b111111, 6'b000111, 6'b111001, 6'b111000, 6'b111110, 6'b000111, 6'b110100, 6'b110110, 6'b001000, 6'b111001, 6'b111000, 6'b001001, 6'b110111, 6'b111101, 6'b001011};
      end
   60: begin
        dout = {6'b000111, 6'b111001, 6'b111000, 6'b111000, 6'b111000, 6'b001010, 6'b000001, 6'b001010, 6'b000111, 6'b111110, 6'b110101, 6'b000011, 6'b111100, 6'b110111, 6'b001010, 6'b001001, 6'b000111, 6'b000101, 6'b001000, 6'b110111, 6'b000110, 6'b001110, 6'b110101, 6'b111000, 6'b000111, 6'b000110, 6'b000100, 6'b111010, 6'b000101, 6'b001011, 6'b000011, 6'b001000};
      end
   61: begin
        dout = {6'b110101, 6'b001010, 6'b110111, 6'b110101, 6'b001000, 6'b001011, 6'b111001, 6'b111101, 6'b000011, 6'b111001, 6'b110111, 6'b111010, 6'b000001, 6'b000101, 6'b010000, 6'b111000, 6'b001000, 6'b111000, 6'b110110, 6'b000010, 6'b001000, 6'b110110, 6'b110110, 6'b111001, 6'b110101, 6'b111100, 6'b000100, 6'b110100, 6'b111001, 6'b001011, 6'b000111, 6'b001001};
      end
   62: begin
        dout = {6'b111101, 6'b110111, 6'b110111, 6'b001001, 6'b001001, 6'b000101, 6'b110111, 6'b000100, 6'b000000, 6'b001110, 6'b001000, 6'b000111, 6'b000010, 6'b111010, 6'b001001, 6'b000101, 6'b000101, 6'b111111, 6'b001001, 6'b110111, 6'b111101, 6'b110101, 6'b111001, 6'b000110, 6'b110110, 6'b101111, 6'b001101, 6'b001000, 6'b110111, 6'b001000, 6'b110011, 6'b111010};
      end
   63: begin
        dout = {6'b110010, 6'b111000, 6'b111101, 6'b001110, 6'b110110, 6'b001000, 6'b001001, 6'b001011, 6'b110101, 6'b000010, 6'b110100, 6'b111000, 6'b111001, 6'b110100, 6'b001001, 6'b110100, 6'b110011, 6'b110110, 6'b001001, 6'b111010, 6'b111010, 6'b110100, 6'b000110, 6'b001001, 6'b001001, 6'b110111, 6'b000111, 6'b111110, 6'b111000, 6'b111101, 6'b111011, 6'b110110};
      end
   64: begin
        dout = {6'b111001, 6'b000100, 6'b000110, 6'b001001, 6'b110000, 6'b110110, 6'b110110, 6'b000010, 6'b111000, 6'b001010, 6'b000100, 6'b001001, 6'b001001, 6'b111010, 6'b001000, 6'b000100, 6'b111001, 6'b000010, 6'b111000, 6'b111111, 6'b000100, 6'b110101, 6'b111000, 6'b110001, 6'b000111, 6'b001000, 6'b111011, 6'b111010, 6'b000100, 6'b000101, 6'b111100, 6'b110110};
      end
   65: begin
        dout = {6'b110110, 6'b110111, 6'b001000, 6'b001000, 6'b001101, 6'b000111, 6'b001011, 6'b111110, 6'b000001, 6'b111000, 6'b001000, 6'b110001, 6'b001000, 6'b110100, 6'b001001, 6'b000110, 6'b111010, 6'b001000, 6'b111001, 6'b001000, 6'b001000, 6'b000110, 6'b101110, 6'b001000, 6'b111001, 6'b111010, 6'b110111, 6'b110110, 6'b001100, 6'b001110, 6'b001001, 6'b000100};
      end
   66: begin
        dout = {6'b111010, 6'b111001, 6'b000100, 6'b110111, 6'b111000, 6'b001000, 6'b110001, 6'b110110, 6'b001110, 6'b001100, 6'b111010, 6'b111001, 6'b001001, 6'b001010, 6'b000011, 6'b111001, 6'b101111, 6'b010001, 6'b110011, 6'b111000, 6'b000100, 6'b111001, 6'b001000, 6'b110100, 6'b110110, 6'b111100, 6'b001010, 6'b000010, 6'b001000, 6'b111000, 6'b110110, 6'b111010};
      end
   67: begin
        dout = {6'b000110, 6'b001010, 6'b000101, 6'b001110, 6'b001111, 6'b110110, 6'b001011, 6'b110111, 6'b001000, 6'b110111, 6'b110011, 6'b000011, 6'b001000, 6'b001000, 6'b110111, 6'b110000, 6'b110011, 6'b110100, 6'b111001, 6'b111000, 6'b001000, 6'b000100, 6'b000110, 6'b111010, 6'b111001, 6'b111000, 6'b110110, 6'b000110, 6'b111001, 6'b111011, 6'b110100, 6'b001110};
      end
   68: begin
        dout = {6'b001100, 6'b001011, 6'b111011, 6'b111010, 6'b000100, 6'b001011, 6'b000111, 6'b000110, 6'b110000, 6'b000101, 6'b111000, 6'b001010, 6'b111100, 6'b000001, 6'b001010, 6'b001100, 6'b001111, 6'b110111, 6'b000101, 6'b001011, 6'b101111, 6'b110010, 6'b000110, 6'b000111, 6'b000110, 6'b111000, 6'b111010, 6'b001000, 6'b001000, 6'b001001, 6'b001101, 6'b110101};
      end
   69: begin
        dout = {6'b111001, 6'b000100, 6'b111001, 6'b110101, 6'b110010, 6'b110100, 6'b111001, 6'b000100, 6'b001001, 6'b001011, 6'b000111, 6'b111101, 6'b111100, 6'b000110, 6'b111011, 6'b110011, 6'b111110, 6'b110110, 6'b111000, 6'b111011, 6'b000001, 6'b001001, 6'b110110, 6'b110000, 6'b110110, 6'b000001, 6'b010000, 6'b110110, 6'b000100, 6'b111000, 6'b111011, 6'b110011};
      end
   70: begin
        dout = {6'b110011, 6'b111101, 6'b110101, 6'b110110, 6'b110100, 6'b111001, 6'b110111, 6'b111010, 6'b110101, 6'b000010, 6'b110011, 6'b000111, 6'b001110, 6'b110101, 6'b111100, 6'b111001, 6'b001001, 6'b110110, 6'b000100, 6'b111001, 6'b110101, 6'b111100, 6'b111001, 6'b000110, 6'b000111, 6'b111110, 6'b000000, 6'b110101, 6'b001101, 6'b110001, 6'b001001, 6'b111000};
      end
   71: begin
        dout = {6'b000010, 6'b110111, 6'b000101, 6'b000110, 6'b000011, 6'b111000, 6'b000110, 6'b000100, 6'b111011, 6'b110101, 6'b001010, 6'b001101, 6'b010000, 6'b000001, 6'b001010, 6'b111110, 6'b000101, 6'b110001, 6'b101101, 6'b111110, 6'b010001, 6'b001100, 6'b000100, 6'b111001, 6'b001011, 6'b111110, 6'b000110, 6'b110101, 6'b001100, 6'b000111, 6'b000001, 6'b001000};
      end
   72: begin
        dout = {6'b111011, 6'b001001, 6'b111010, 6'b110110, 6'b000110, 6'b111011, 6'b001000, 6'b111001, 6'b001010, 6'b111000, 6'b111100, 6'b000001, 6'b110011, 6'b111110, 6'b111001, 6'b000110, 6'b000110, 6'b110000, 6'b000110, 6'b110111, 6'b000110, 6'b110011, 6'b111100, 6'b001011, 6'b110110, 6'b111000, 6'b111001, 6'b110100, 6'b000100, 6'b111010, 6'b001101, 6'b111111};
      end
   73: begin
        dout = {6'b111000, 6'b110000, 6'b001010, 6'b110001, 6'b001000, 6'b110000, 6'b110101, 6'b111011, 6'b000110, 6'b110000, 6'b000100, 6'b010000, 6'b000100, 6'b110001, 6'b001010, 6'b101111, 6'b001000, 6'b111010, 6'b111010, 6'b001001, 6'b110101, 6'b001010, 6'b001000, 6'b111011, 6'b110111, 6'b110111, 6'b000100, 6'b111100, 6'b111100, 6'b111110, 6'b110011, 6'b000101};
      end
   74: begin
        dout = {6'b110111, 6'b110011, 6'b001000, 6'b110101, 6'b110101, 6'b000011, 6'b001110, 6'b001110, 6'b111101, 6'b000101, 6'b001000, 6'b111010, 6'b111000, 6'b110100, 6'b111001, 6'b111010, 6'b000110, 6'b111001, 6'b001111, 6'b111000, 6'b001001, 6'b111110, 6'b111001, 6'b110110, 6'b111111, 6'b001001, 6'b000111, 6'b111000, 6'b001000, 6'b110010, 6'b000111, 6'b001000};
      end
   75: begin
        dout = {6'b001101, 6'b000000, 6'b110111, 6'b001001, 6'b000110, 6'b110111, 6'b000111, 6'b000101, 6'b001001, 6'b111010, 6'b110111, 6'b001010, 6'b001011, 6'b111001, 6'b001110, 6'b111011, 6'b001011, 6'b111101, 6'b001010, 6'b001010, 6'b111000, 6'b110110, 6'b001011, 6'b110010, 6'b110101, 6'b110000, 6'b101110, 6'b111001, 6'b110011, 6'b000111, 6'b001101, 6'b110111};
      end
   76: begin
        dout = {6'b111001, 6'b001101, 6'b000110, 6'b000100, 6'b000001, 6'b001011, 6'b000101, 6'b001010, 6'b111001, 6'b111001, 6'b000110, 6'b001011, 6'b101111, 6'b111001, 6'b110100, 6'b111110, 6'b111010, 6'b000001, 6'b000101, 6'b001101, 6'b111001, 6'b110010, 6'b111111, 6'b110011, 6'b101111, 6'b110101, 6'b111110, 6'b000111, 6'b001010, 6'b001000, 6'b110101, 6'b110111};
      end
   77: begin
        dout = {6'b111111, 6'b000110, 6'b110110, 6'b111000, 6'b111110, 6'b001001, 6'b001111, 6'b111000, 6'b111001, 6'b001100, 6'b110110, 6'b000110, 6'b111010, 6'b110010, 6'b001111, 6'b110110, 6'b110111, 6'b111111, 6'b001011, 6'b111010, 6'b110100, 6'b000101, 6'b001001, 6'b000110, 6'b001001, 6'b110111, 6'b001110, 6'b111100, 6'b110011, 6'b111000, 6'b110110, 6'b110111};
      end
   78: begin
        dout = {6'b001000, 6'b111000, 6'b110111, 6'b111010, 6'b110100, 6'b111010, 6'b000100, 6'b111010, 6'b001000, 6'b110100, 6'b110100, 6'b001000, 6'b111001, 6'b111001, 6'b001100, 6'b111001, 6'b110110, 6'b111011, 6'b110010, 6'b110110, 6'b111100, 6'b111100, 6'b001100, 6'b110111, 6'b111000, 6'b001010, 6'b000110, 6'b001001, 6'b000111, 6'b111001, 6'b001111, 6'b111001};
      end
   79: begin
        dout = {6'b001100, 6'b110001, 6'b111101, 6'b001000, 6'b111101, 6'b000101, 6'b001010, 6'b000100, 6'b001010, 6'b001101, 6'b000001, 6'b110101, 6'b001001, 6'b001010, 6'b110100, 6'b110110, 6'b110100, 6'b001010, 6'b000100, 6'b110000, 6'b010001, 6'b111011, 6'b000100, 6'b111001, 6'b110111, 6'b111000, 6'b000101, 6'b000100, 6'b111001, 6'b001010, 6'b111000, 6'b001000};
      end
   80: begin
        dout = {6'b000100, 6'b111100, 6'b000100, 6'b000100, 6'b111000, 6'b001010, 6'b001001, 6'b001011, 6'b111001, 6'b000100, 6'b111100, 6'b000110, 6'b001000, 6'b111000, 6'b001001, 6'b111001, 6'b001100, 6'b010110, 6'b110001, 6'b001001, 6'b111110, 6'b110100, 6'b111110, 6'b000101, 6'b110101, 6'b000101, 6'b110011, 6'b000111, 6'b001011, 6'b111011, 6'b000110, 6'b111000};
      end
   81: begin
        dout = {6'b001100, 6'b001000, 6'b000101, 6'b110111, 6'b111001, 6'b110111, 6'b001101, 6'b000011, 6'b000110, 6'b000110, 6'b111011, 6'b110110, 6'b000001, 6'b111001, 6'b000110, 6'b111000, 6'b110010, 6'b000110, 6'b110111, 6'b110101, 6'b110111, 6'b000111, 6'b110110, 6'b111001, 6'b111001, 6'b110111, 6'b111010, 6'b000001, 6'b110010, 6'b000111, 6'b110111, 6'b001001};
      end
   82: begin
        dout = {6'b000110, 6'b110001, 6'b000011, 6'b110011, 6'b111000, 6'b111000, 6'b111001, 6'b111001, 6'b000101, 6'b110111, 6'b001010, 6'b001010, 6'b001010, 6'b001000, 6'b000111, 6'b111100, 6'b010000, 6'b110110, 6'b001011, 6'b111011, 6'b000100, 6'b000011, 6'b111000, 6'b000110, 6'b001010, 6'b000101, 6'b111111, 6'b000100, 6'b001101, 6'b001000, 6'b000101, 6'b110110};
      end
   83: begin
        dout = {6'b000010, 6'b000110, 6'b110100, 6'b111001, 6'b000101, 6'b001111, 6'b000100, 6'b111001, 6'b110100, 6'b110101, 6'b110001, 6'b001001, 6'b110111, 6'b101101, 6'b110100, 6'b000011, 6'b000101, 6'b111100, 6'b110001, 6'b111110, 6'b000001, 6'b111100, 6'b110111, 6'b000111, 6'b111000, 6'b111011, 6'b111001, 6'b111001, 6'b001010, 6'b000101, 6'b110101, 6'b111111};
      end
   84: begin
        dout = {6'b111101, 6'b001101, 6'b111011, 6'b110111, 6'b000100, 6'b111001, 6'b001010, 6'b001111, 6'b001000, 6'b001101, 6'b001011, 6'b000101, 6'b111100, 6'b110100, 6'b000100, 6'b110111, 6'b001010, 6'b000100, 6'b110111, 6'b111101, 6'b111010, 6'b110101, 6'b001000, 6'b001101, 6'b001010, 6'b111101, 6'b111000, 6'b110100, 6'b110110, 6'b111010, 6'b001010, 6'b110100};
      end
   85: begin
        dout = {6'b111010, 6'b001011, 6'b111001, 6'b111110, 6'b110110, 6'b000101, 6'b110111, 6'b111000, 6'b000101, 6'b111001, 6'b101111, 6'b000110, 6'b001000, 6'b111010, 6'b000100, 6'b001101, 6'b001001, 6'b111011, 6'b110110, 6'b001000, 6'b101100, 6'b001100, 6'b110111, 6'b111011, 6'b110101, 6'b111000, 6'b110111, 6'b000100, 6'b000110, 6'b111001, 6'b111001, 6'b110111};
      end
   86: begin
        dout = {6'b000100, 6'b110111, 6'b001000, 6'b000010, 6'b000100, 6'b110011, 6'b111001, 6'b000101, 6'b000101, 6'b000011, 6'b110101, 6'b111010, 6'b001000, 6'b111101, 6'b001001, 6'b110111, 6'b000101, 6'b000111, 6'b110101, 6'b000010, 6'b111010, 6'b001101, 6'b000001, 6'b000110, 6'b001100, 6'b010000, 6'b111000, 6'b110101, 6'b000101, 6'b001000, 6'b001010, 6'b110010};
      end
   87: begin
        dout = {6'b000100, 6'b111001, 6'b110110, 6'b001000, 6'b000101, 6'b001010, 6'b111001, 6'b110001, 6'b001000, 6'b000110, 6'b000110, 6'b111101, 6'b111000, 6'b110010, 6'b111101, 6'b111010, 6'b001101, 6'b111100, 6'b110111, 6'b001101, 6'b010000, 6'b000001, 6'b110110, 6'b001001, 6'b110010, 6'b110101, 6'b000111, 6'b110011, 6'b000100, 6'b000100, 6'b000110, 6'b001001};
      end
   88: begin
        dout = {6'b111100, 6'b110001, 6'b000010, 6'b000101, 6'b000100, 6'b111111, 6'b110110, 6'b110110, 6'b000100, 6'b111010, 6'b111000, 6'b111110, 6'b111110, 6'b001010, 6'b000101, 6'b000010, 6'b000101, 6'b111001, 6'b110101, 6'b000110, 6'b000001, 6'b001010, 6'b110101, 6'b111001, 6'b111000, 6'b111000, 6'b001111, 6'b001100, 6'b001010, 6'b001000, 6'b001101, 6'b111001};
      end
   89: begin
        dout = {6'b110101, 6'b000111, 6'b111010, 6'b000010, 6'b001110, 6'b001100, 6'b001100, 6'b001000, 6'b111010, 6'b001010, 6'b001011, 6'b110100, 6'b111001, 6'b111001, 6'b001000, 6'b000011, 6'b001001, 6'b000010, 6'b110111, 6'b000100, 6'b000101, 6'b000110, 6'b111001, 6'b110111, 6'b111101, 6'b001000, 6'b110110, 6'b110010, 6'b001101, 6'b000111, 6'b110111, 6'b110111};
      end
   90: begin
        dout = {6'b110011, 6'b110111, 6'b001000, 6'b111000, 6'b001001, 6'b000010, 6'b111010, 6'b000100, 6'b000110, 6'b000100, 6'b111010, 6'b110110, 6'b111001, 6'b110101, 6'b110011, 6'b000110, 6'b000100, 6'b110010, 6'b001001, 6'b001010, 6'b001110, 6'b001001, 6'b000010, 6'b000010, 6'b110110, 6'b000111, 6'b000111, 6'b110110, 6'b110110, 6'b001111, 6'b110111, 6'b001111};
      end
   91: begin
        dout = {6'b111101, 6'b000110, 6'b000111, 6'b001101, 6'b001000, 6'b000100, 6'b110111, 6'b000111, 6'b111010, 6'b111001, 6'b111110, 6'b110111, 6'b001100, 6'b001110, 6'b000111, 6'b111011, 6'b110101, 6'b110100, 6'b001100, 6'b110110, 6'b000111, 6'b001010, 6'b110111, 6'b001010, 6'b000101, 6'b111101, 6'b111110, 6'b110100, 6'b111010, 6'b000101, 6'b110101, 6'b001011};
      end
   92: begin
        dout = {6'b110111, 6'b001000, 6'b110111, 6'b110100, 6'b001100, 6'b000110, 6'b000001, 6'b000110, 6'b001011, 6'b000111, 6'b110110, 6'b110011, 6'b111001, 6'b000110, 6'b000011, 6'b110000, 6'b110101, 6'b000110, 6'b110111, 6'b110110, 6'b110010, 6'b110110, 6'b000100, 6'b000110, 6'b000010, 6'b111000, 6'b000111, 6'b110010, 6'b001101, 6'b001000, 6'b000110, 6'b110101};
      end
   93: begin
        dout = {6'b111010, 6'b001110, 6'b111101, 6'b001001, 6'b001100, 6'b000111, 6'b000110, 6'b000100, 6'b000011, 6'b001100, 6'b110110, 6'b111010, 6'b000100, 6'b001011, 6'b110110, 6'b110010, 6'b111010, 6'b111101, 6'b000100, 6'b001110, 6'b000111, 6'b111111, 6'b110111, 6'b111001, 6'b110101, 6'b000001, 6'b001101, 6'b000110, 6'b110111, 6'b000011, 6'b110100, 6'b000101};
      end
   94: begin
        dout = {6'b001001, 6'b110110, 6'b000101, 6'b000101, 6'b110111, 6'b111101, 6'b110110, 6'b110110, 6'b000110, 6'b000000, 6'b110101, 6'b111011, 6'b110111, 6'b111000, 6'b111001, 6'b000001, 6'b110001, 6'b111010, 6'b111000, 6'b111001, 6'b110111, 6'b000101, 6'b111110, 6'b000011, 6'b111100, 6'b000110, 6'b111001, 6'b000100, 6'b000010, 6'b000110, 6'b111010, 6'b111000};
      end
   95: begin
        dout = {6'b110111, 6'b001010, 6'b000001, 6'b110111, 6'b001000, 6'b000100, 6'b000000, 6'b001111, 6'b111000, 6'b000101, 6'b000111, 6'b111011, 6'b110111, 6'b110110, 6'b110110, 6'b001000, 6'b000111, 6'b000111, 6'b001010, 6'b000101, 6'b111010, 6'b111001, 6'b111001, 6'b111111, 6'b000010, 6'b000101, 6'b001011, 6'b111001, 6'b111000, 6'b111011, 6'b111001, 6'b111001};
      end
   96: begin
        dout = {6'b111111, 6'b110000, 6'b110010, 6'b000111, 6'b111001, 6'b000011, 6'b110101, 6'b001011, 6'b001001, 6'b111100, 6'b001010, 6'b111010, 6'b001100, 6'b111010, 6'b000110, 6'b000101, 6'b001100, 6'b001100, 6'b111101, 6'b111010, 6'b001010, 6'b001101, 6'b000110, 6'b001001, 6'b001111, 6'b111001, 6'b111110, 6'b000100, 6'b000110, 6'b110100, 6'b111010, 6'b111101};
      end
   97: begin
        dout = {6'b111101, 6'b111000, 6'b001010, 6'b000100, 6'b111110, 6'b101111, 6'b000111, 6'b110100, 6'b001101, 6'b110100, 6'b110111, 6'b110010, 6'b001100, 6'b001001, 6'b001001, 6'b110011, 6'b110010, 6'b110110, 6'b110111, 6'b110110, 6'b000110, 6'b110011, 6'b111011, 6'b110110, 6'b111101, 6'b000110, 6'b111000, 6'b000100, 6'b110000, 6'b001011, 6'b110111, 6'b111010};
      end
   98: begin
        dout = {6'b111010, 6'b000011, 6'b001100, 6'b001011, 6'b111011, 6'b000111, 6'b111010, 6'b110101, 6'b001111, 6'b001001, 6'b000100, 6'b001000, 6'b110110, 6'b110110, 6'b000001, 6'b111000, 6'b111010, 6'b000111, 6'b111000, 6'b110011, 6'b000110, 6'b111000, 6'b111010, 6'b000110, 6'b001011, 6'b111010, 6'b110110, 6'b111000, 6'b000100, 6'b111110, 6'b111001, 6'b000100};
      end
   99: begin
        dout = {6'b001100, 6'b001001, 6'b001001, 6'b001010, 6'b001111, 6'b000110, 6'b110010, 6'b000101, 6'b001000, 6'b001100, 6'b111010, 6'b110111, 6'b111110, 6'b000101, 6'b111100, 6'b110101, 6'b110111, 6'b111010, 6'b110110, 6'b110111, 6'b110100, 6'b111001, 6'b110101, 6'b110010, 6'b001101, 6'b111100, 6'b001011, 6'b111010, 6'b110011, 6'b110001, 6'b000010, 6'b001100};
      end
   100: begin
        dout = {6'b111011, 6'b001011, 6'b001110, 6'b000101, 6'b111001, 6'b001010, 6'b110010, 6'b110101, 6'b111011, 6'b001010, 6'b110110, 6'b000010, 6'b110111, 6'b110011, 6'b111101, 6'b111011, 6'b001000, 6'b000010, 6'b000000, 6'b001001, 6'b110100, 6'b000110, 6'b000001, 6'b001001, 6'b000101, 6'b000111, 6'b110111, 6'b001100, 6'b110100, 6'b111000, 6'b111110, 6'b001101};
      end
   101: begin
        dout = {6'b111100, 6'b110011, 6'b000100, 6'b000011, 6'b111010, 6'b110110, 6'b000010, 6'b001011, 6'b001011, 6'b001010, 6'b111000, 6'b001010, 6'b110110, 6'b000111, 6'b101111, 6'b111100, 6'b110011, 6'b110100, 6'b000101, 6'b001100, 6'b001100, 6'b001000, 6'b000110, 6'b110100, 6'b110101, 6'b111110, 6'b110110, 6'b000011, 6'b000100, 6'b110011, 6'b111010, 6'b001011};
      end
   102: begin
        dout = {6'b000011, 6'b110111, 6'b110111, 6'b001111, 6'b000100, 6'b111100, 6'b110010, 6'b110011, 6'b001001, 6'b110011, 6'b000011, 6'b001000, 6'b000011, 6'b000100, 6'b111100, 6'b110110, 6'b000100, 6'b110110, 6'b111001, 6'b000011, 6'b110100, 6'b111000, 6'b110011, 6'b000101, 6'b110111, 6'b110111, 6'b010001, 6'b000101, 6'b000000, 6'b110001, 6'b000011, 6'b111010};
      end
   103: begin
        dout = {6'b001001, 6'b111000, 6'b000011, 6'b000110, 6'b000001, 6'b000100, 6'b111001, 6'b111010, 6'b000100, 6'b001010, 6'b110001, 6'b110011, 6'b000001, 6'b001001, 6'b111000, 6'b111001, 6'b110101, 6'b110101, 6'b111010, 6'b111011, 6'b000111, 6'b001010, 6'b000111, 6'b110010, 6'b000011, 6'b111010, 6'b111010, 6'b000100, 6'b111001, 6'b000001, 6'b001000, 6'b001010};
      end
   104: begin
        dout = {6'b000101, 6'b001100, 6'b110011, 6'b000100, 6'b000010, 6'b111000, 6'b110111, 6'b000011, 6'b001101, 6'b001011, 6'b000110, 6'b000100, 6'b110011, 6'b000111, 6'b111001, 6'b110110, 6'b110100, 6'b110101, 6'b110011, 6'b111000, 6'b000101, 6'b110101, 6'b110010, 6'b110010, 6'b000101, 6'b110001, 6'b001001, 6'b000100, 6'b110111, 6'b001100, 6'b001011, 6'b001100};
      end
   105: begin
        dout = {6'b000111, 6'b111001, 6'b001000, 6'b111100, 6'b000111, 6'b000100, 6'b001010, 6'b000101, 6'b110101, 6'b111110, 6'b110110, 6'b000010, 6'b001011, 6'b111010, 6'b001000, 6'b111100, 6'b110111, 6'b110011, 6'b000111, 6'b000110, 6'b000101, 6'b000001, 6'b001010, 6'b000111, 6'b000110, 6'b111111, 6'b111011, 6'b111100, 6'b001111, 6'b111001, 6'b000011, 6'b111010};
      end
   106: begin
        dout = {6'b000011, 6'b001011, 6'b110111, 6'b001000, 6'b001100, 6'b000111, 6'b000111, 6'b111000, 6'b001010, 6'b000100, 6'b111010, 6'b111011, 6'b110100, 6'b110100, 6'b000010, 6'b000001, 6'b110111, 6'b001010, 6'b001000, 6'b001010, 6'b000011, 6'b001110, 6'b110101, 6'b110100, 6'b001000, 6'b111101, 6'b111001, 6'b000010, 6'b000001, 6'b110100, 6'b010000, 6'b111100};
      end
   107: begin
        dout = {6'b000111, 6'b110110, 6'b111001, 6'b001010, 6'b001001, 6'b110101, 6'b001010, 6'b001010, 6'b111100, 6'b000010, 6'b000111, 6'b110101, 6'b110110, 6'b111001, 6'b110010, 6'b000100, 6'b010001, 6'b111000, 6'b111011, 6'b001001, 6'b010000, 6'b001100, 6'b110100, 6'b110101, 6'b110101, 6'b000100, 6'b111001, 6'b110001, 6'b001000, 6'b000010, 6'b000111, 6'b110001};
      end
   108: begin
        dout = {6'b111010, 6'b111110, 6'b110101, 6'b000010, 6'b110100, 6'b000111, 6'b001010, 6'b000111, 6'b111110, 6'b110111, 6'b000010, 6'b000010, 6'b001000, 6'b111101, 6'b001000, 6'b001000, 6'b000011, 6'b110100, 6'b110111, 6'b000010, 6'b000001, 6'b111000, 6'b001000, 6'b001000, 6'b110100, 6'b111000, 6'b110111, 6'b000110, 6'b110101, 6'b111010, 6'b110111, 6'b000110};
      end
   109: begin
        dout = {6'b001001, 6'b111010, 6'b000110, 6'b001101, 6'b111000, 6'b001010, 6'b001010, 6'b001000, 6'b111100, 6'b001101, 6'b000011, 6'b111100, 6'b001011, 6'b001010, 6'b111110, 6'b000110, 6'b111001, 6'b110111, 6'b110100, 6'b110111, 6'b111011, 6'b111110, 6'b000110, 6'b101111, 6'b110110, 6'b111011, 6'b110101, 6'b000111, 6'b000100, 6'b000111, 6'b111000, 6'b111000};
      end
   110: begin
        dout = {6'b000000, 6'b001001, 6'b110100, 6'b111000, 6'b111101, 6'b000001, 6'b001010, 6'b111001, 6'b001010, 6'b001001, 6'b000101, 6'b110111, 6'b001000, 6'b010000, 6'b111001, 6'b111010, 6'b000101, 6'b000011, 6'b111001, 6'b000101, 6'b111001, 6'b001101, 6'b110110, 6'b001001, 6'b001001, 6'b010000, 6'b110100, 6'b001100, 6'b000101, 6'b111101, 6'b111010, 6'b000110};
      end
   111: begin
        dout = {6'b111011, 6'b111000, 6'b110110, 6'b001010, 6'b110110, 6'b001010, 6'b110111, 6'b111001, 6'b000011, 6'b001001, 6'b001001, 6'b111011, 6'b001100, 6'b111010, 6'b000111, 6'b111000, 6'b101101, 6'b001010, 6'b000111, 6'b110111, 6'b000111, 6'b110101, 6'b001110, 6'b000110, 6'b001101, 6'b001111, 6'b110111, 6'b001011, 6'b110110, 6'b000100, 6'b111000, 6'b000100};
      end
   112: begin
        dout = {6'b111001, 6'b001000, 6'b001010, 6'b000100, 6'b110110, 6'b001000, 6'b001000, 6'b001011, 6'b110110, 6'b110110, 6'b001001, 6'b001010, 6'b000100, 6'b000000, 6'b001100, 6'b111100, 6'b000010, 6'b000100, 6'b111001, 6'b000111, 6'b110111, 6'b001001, 6'b001101, 6'b000111, 6'b111000, 6'b000100, 6'b111101, 6'b110101, 6'b001110, 6'b111010, 6'b110101, 6'b111001};
      end
   113: begin
        dout = {6'b111111, 6'b111010, 6'b111001, 6'b110010, 6'b001001, 6'b000110, 6'b001100, 6'b110001, 6'b110011, 6'b001100, 6'b001111, 6'b000111, 6'b001100, 6'b111110, 6'b111001, 6'b111001, 6'b000101, 6'b000011, 6'b111000, 6'b001000, 6'b000111, 6'b001000, 6'b001011, 6'b110111, 6'b111001, 6'b000100, 6'b110011, 6'b111001, 6'b111000, 6'b111001, 6'b111000, 6'b111000};
      end
   114: begin
        dout = {6'b000011, 6'b111010, 6'b111101, 6'b110110, 6'b111101, 6'b110100, 6'b001110, 6'b111011, 6'b111000, 6'b000010, 6'b110111, 6'b000100, 6'b000100, 6'b111000, 6'b111001, 6'b111100, 6'b001001, 6'b111011, 6'b000110, 6'b111111, 6'b001000, 6'b000110, 6'b111000, 6'b110001, 6'b110110, 6'b001110, 6'b001000, 6'b111101, 6'b001000, 6'b111000, 6'b111000, 6'b110110};
      end
   115: begin
        dout = {6'b000101, 6'b000110, 6'b001000, 6'b001101, 6'b110010, 6'b111110, 6'b111010, 6'b000100, 6'b001001, 6'b110110, 6'b001001, 6'b110010, 6'b001100, 6'b000100, 6'b000101, 6'b110010, 6'b001011, 6'b001001, 6'b110000, 6'b000011, 6'b001010, 6'b110100, 6'b000101, 6'b000101, 6'b110111, 6'b110101, 6'b000111, 6'b111000, 6'b110011, 6'b111011, 6'b110010, 6'b110110};
      end
   116: begin
        dout = {6'b111101, 6'b111001, 6'b111011, 6'b111000, 6'b110110, 6'b110110, 6'b000110, 6'b111011, 6'b001110, 6'b111001, 6'b110111, 6'b000110, 6'b000110, 6'b000110, 6'b000111, 6'b110110, 6'b000110, 6'b111000, 6'b000101, 6'b001000, 6'b110110, 6'b111011, 6'b000111, 6'b000110, 6'b000101, 6'b110011, 6'b110100, 6'b000111, 6'b111010, 6'b000101, 6'b000011, 6'b000101};
      end
   117: begin
        dout = {6'b111100, 6'b110011, 6'b110110, 6'b001001, 6'b001011, 6'b001101, 6'b000110, 6'b111101, 6'b110011, 6'b001011, 6'b001111, 6'b111001, 6'b000111, 6'b000011, 6'b001100, 6'b111101, 6'b111000, 6'b000100, 6'b000111, 6'b001100, 6'b110110, 6'b001010, 6'b110111, 6'b001111, 6'b001001, 6'b001110, 6'b000000, 6'b111101, 6'b111011, 6'b000110, 6'b110011, 6'b001011};
      end
   118: begin
        dout = {6'b110111, 6'b000100, 6'b001001, 6'b111110, 6'b000111, 6'b111010, 6'b110110, 6'b110101, 6'b111101, 6'b110100, 6'b110111, 6'b000000, 6'b110110, 6'b111000, 6'b001010, 6'b110110, 6'b111000, 6'b111001, 6'b101111, 6'b001010, 6'b111110, 6'b111000, 6'b000110, 6'b001101, 6'b001001, 6'b110010, 6'b110111, 6'b001010, 6'b110101, 6'b110110, 6'b001000, 6'b000111};
      end
   119: begin
        dout = {6'b110011, 6'b000001, 6'b001001, 6'b111000, 6'b110111, 6'b111111, 6'b110111, 6'b001010, 6'b001001, 6'b111000, 6'b110101, 6'b110110, 6'b000110, 6'b001111, 6'b001000, 6'b000110, 6'b110100, 6'b001100, 6'b111100, 6'b001110, 6'b111011, 6'b110111, 6'b110111, 6'b001010, 6'b000101, 6'b111000, 6'b001001, 6'b111001, 6'b000010, 6'b110111, 6'b001000, 6'b001100};
      end
   120: begin
        dout = {6'b001010, 6'b001000, 6'b001101, 6'b110111, 6'b110011, 6'b110111, 6'b001001, 6'b101110, 6'b111010, 6'b001000, 6'b111000, 6'b110101, 6'b110111, 6'b001010, 6'b110111, 6'b110111, 6'b110101, 6'b000110, 6'b000101, 6'b001101, 6'b001000, 6'b111010, 6'b111111, 6'b111001, 6'b000101, 6'b111000, 6'b111111, 6'b000100, 6'b000100, 6'b110110, 6'b111101, 6'b111011};
      end
   121: begin
        dout = {6'b000100, 6'b110010, 6'b110110, 6'b000100, 6'b110100, 6'b000011, 6'b000101, 6'b110011, 6'b000101, 6'b110110, 6'b111010, 6'b001000, 6'b111010, 6'b110100, 6'b110101, 6'b000011, 6'b110111, 6'b110110, 6'b000101, 6'b000010, 6'b111101, 6'b001101, 6'b111110, 6'b111101, 6'b110111, 6'b001001, 6'b111000, 6'b111010, 6'b110101, 6'b111010, 6'b110100, 6'b111100};
      end
   122: begin
        dout = {6'b111001, 6'b000001, 6'b000000, 6'b111011, 6'b001000, 6'b111001, 6'b111100, 6'b111011, 6'b111010, 6'b110010, 6'b111010, 6'b110101, 6'b111001, 6'b000101, 6'b111010, 6'b110110, 6'b000011, 6'b001001, 6'b111011, 6'b001010, 6'b001001, 6'b110111, 6'b000110, 6'b111000, 6'b000101, 6'b001010, 6'b000000, 6'b000111, 6'b111110, 6'b110110, 6'b000110, 6'b110010};
      end
   123: begin
        dout = {6'b000101, 6'b000111, 6'b001010, 6'b111100, 6'b111000, 6'b111000, 6'b111100, 6'b111001, 6'b110101, 6'b110011, 6'b110100, 6'b001010, 6'b001001, 6'b110010, 6'b000101, 6'b000110, 6'b111001, 6'b111011, 6'b001101, 6'b000101, 6'b001011, 6'b000111, 6'b000101, 6'b110101, 6'b001001, 6'b110101, 6'b111011, 6'b110010, 6'b110001, 6'b001000, 6'b000110, 6'b000011};
      end
   124: begin
        dout = {6'b000110, 6'b110111, 6'b001011, 6'b110101, 6'b001101, 6'b111100, 6'b111100, 6'b111010, 6'b010001, 6'b001101, 6'b000100, 6'b000101, 6'b111001, 6'b110111, 6'b110011, 6'b001010, 6'b110111, 6'b110101, 6'b110110, 6'b110111, 6'b111000, 6'b000101, 6'b000111, 6'b101110, 6'b001011, 6'b111001, 6'b111100, 6'b110111, 6'b000100, 6'b001010, 6'b111010, 6'b110111};
      end
   125: begin
        dout = {6'b000110, 6'b111101, 6'b111001, 6'b111000, 6'b111000, 6'b001100, 6'b111001, 6'b110100, 6'b110011, 6'b111000, 6'b110111, 6'b111010, 6'b111100, 6'b001010, 6'b001000, 6'b111010, 6'b001110, 6'b111100, 6'b001000, 6'b001101, 6'b111001, 6'b001001, 6'b010000, 6'b111001, 6'b001010, 6'b001010, 6'b000111, 6'b001011, 6'b110100, 6'b111010, 6'b000100, 6'b001100};
      end
   126: begin
        dout = {6'b110110, 6'b101110, 6'b000101, 6'b000111, 6'b001110, 6'b001010, 6'b000110, 6'b001010, 6'b111101, 6'b000100, 6'b000100, 6'b001010, 6'b110111, 6'b000111, 6'b111011, 6'b000011, 6'b111010, 6'b111011, 6'b000111, 6'b000101, 6'b110110, 6'b110110, 6'b111000, 6'b001101, 6'b001110, 6'b001001, 6'b001000, 6'b001010, 6'b001001, 6'b000101, 6'b110101, 6'b110110};
      end
   127: begin
        dout = {6'b001001, 6'b101111, 6'b111000, 6'b000110, 6'b000010, 6'b111110, 6'b111001, 6'b101101, 6'b110011, 6'b110110, 6'b111000, 6'b111010, 6'b110110, 6'b001001, 6'b000110, 6'b111110, 6'b110110, 6'b110110, 6'b000011, 6'b000110, 6'b110011, 6'b110111, 6'b110100, 6'b110110, 6'b111100, 6'b000110, 6'b001010, 6'b000110, 6'b000100, 6'b110011, 6'b000110, 6'b111000};
      end
   128: begin
        dout = {6'b000101, 6'b111000, 6'b110100, 6'b001001, 6'b110111, 6'b110100, 6'b001000, 6'b001010, 6'b000100, 6'b000111, 6'b001000, 6'b110111, 6'b110100, 6'b111001, 6'b111111, 6'b110111, 6'b111110, 6'b001010, 6'b110101, 6'b001010, 6'b111111, 6'b001011, 6'b001010, 6'b001001, 6'b111010, 6'b110100, 6'b110010, 6'b000010, 6'b111001, 6'b110011, 6'b110111, 6'b001001};
      end
   129: begin
        dout = {6'b110101, 6'b110100, 6'b001000, 6'b001000, 6'b111100, 6'b111100, 6'b001001, 6'b111100, 6'b111010, 6'b000111, 6'b110111, 6'b111110, 6'b000101, 6'b010000, 6'b111011, 6'b000110, 6'b001011, 6'b000111, 6'b110010, 6'b001100, 6'b000011, 6'b001110, 6'b000100, 6'b110101, 6'b000100, 6'b001000, 6'b000110, 6'b110011, 6'b001010, 6'b001001, 6'b000101, 6'b110111};
      end
   130: begin
        dout = {6'b111001, 6'b001100, 6'b000011, 6'b111001, 6'b001000, 6'b111111, 6'b110010, 6'b111000, 6'b000110, 6'b000110, 6'b110111, 6'b110100, 6'b001011, 6'b000111, 6'b001000, 6'b111101, 6'b110110, 6'b000011, 6'b110111, 6'b110011, 6'b111001, 6'b000011, 6'b001011, 6'b001001, 6'b000111, 6'b111111, 6'b111010, 6'b000101, 6'b111101, 6'b001011, 6'b111011, 6'b110011};
      end
   131: begin
        dout = {6'b000101, 6'b101111, 6'b111011, 6'b000110, 6'b000111, 6'b001001, 6'b000010, 6'b000100, 6'b110111, 6'b111100, 6'b110010, 6'b111010, 6'b000100, 6'b111010, 6'b111011, 6'b111010, 6'b001100, 6'b001000, 6'b111010, 6'b001010, 6'b000011, 6'b110101, 6'b111111, 6'b000101, 6'b110010, 6'b001100, 6'b110111, 6'b111001, 6'b110111, 6'b111100, 6'b111100, 6'b110100};
      end
   132: begin
        dout = {6'b000100, 6'b110010, 6'b001100, 6'b111111, 6'b110100, 6'b110110, 6'b111111, 6'b000101, 6'b111011, 6'b111010, 6'b111100, 6'b101110, 6'b111111, 6'b001111, 6'b001101, 6'b111010, 6'b110010, 6'b110101, 6'b110111, 6'b000111, 6'b000001, 6'b001011, 6'b110000, 6'b111000, 6'b111110, 6'b111010, 6'b001001, 6'b111100, 6'b110111, 6'b001011, 6'b111010, 6'b001100};
      end
   133: begin
        dout = {6'b001100, 6'b001010, 6'b111001, 6'b000111, 6'b110101, 6'b000111, 6'b001101, 6'b110111, 6'b111000, 6'b111110, 6'b111000, 6'b001110, 6'b101101, 6'b000111, 6'b110110, 6'b000111, 6'b000101, 6'b111110, 6'b110101, 6'b001101, 6'b110110, 6'b001001, 6'b111010, 6'b001010, 6'b110100, 6'b110111, 6'b110110, 6'b111000, 6'b110111, 6'b000110, 6'b110111, 6'b000100};
      end
   134: begin
        dout = {6'b000010, 6'b111011, 6'b110011, 6'b111010, 6'b000101, 6'b000110, 6'b000101, 6'b001110, 6'b001011, 6'b110111, 6'b110111, 6'b111011, 6'b111001, 6'b001001, 6'b000011, 6'b000001, 6'b000100, 6'b110111, 6'b110100, 6'b111010, 6'b001111, 6'b110110, 6'b001010, 6'b000100, 6'b110110, 6'b001000, 6'b110101, 6'b000111, 6'b010010, 6'b001100, 6'b000110, 6'b111101};
      end
   135: begin
        dout = {6'b110101, 6'b001100, 6'b110101, 6'b000110, 6'b001001, 6'b110001, 6'b110011, 6'b111101, 6'b001000, 6'b000100, 6'b110101, 6'b010001, 6'b001001, 6'b001100, 6'b111001, 6'b111001, 6'b111110, 6'b110111, 6'b000001, 6'b111010, 6'b001000, 6'b001010, 6'b110001, 6'b001100, 6'b111001, 6'b000100, 6'b000010, 6'b111011, 6'b001000, 6'b110100, 6'b110011, 6'b111011};
      end
   136: begin
        dout = {6'b110110, 6'b111100, 6'b001000, 6'b001101, 6'b110101, 6'b001011, 6'b000111, 6'b001001, 6'b001010, 6'b001101, 6'b000111, 6'b110110, 6'b101110, 6'b110100, 6'b000001, 6'b110011, 6'b001000, 6'b001001, 6'b110011, 6'b001000, 6'b000010, 6'b110010, 6'b000101, 6'b110010, 6'b110101, 6'b111010, 6'b111101, 6'b111100, 6'b001001, 6'b000001, 6'b110111, 6'b111000};
      end
   137: begin
        dout = {6'b001001, 6'b110001, 6'b111101, 6'b000101, 6'b111001, 6'b001010, 6'b001001, 6'b001100, 6'b110110, 6'b110100, 6'b001000, 6'b110111, 6'b111001, 6'b000110, 6'b000111, 6'b111011, 6'b110101, 6'b111100, 6'b110110, 6'b110100, 6'b110100, 6'b110100, 6'b000100, 6'b001010, 6'b000001, 6'b000111, 6'b110111, 6'b000001, 6'b110010, 6'b001010, 6'b111001, 6'b001110};
      end
   138: begin
        dout = {6'b001100, 6'b110101, 6'b000111, 6'b000110, 6'b110110, 6'b110111, 6'b110101, 6'b000110, 6'b110010, 6'b110110, 6'b111001, 6'b111101, 6'b000101, 6'b001011, 6'b110110, 6'b110101, 6'b001110, 6'b001001, 6'b111011, 6'b111001, 6'b111011, 6'b000101, 6'b000111, 6'b110011, 6'b111101, 6'b000011, 6'b001100, 6'b110110, 6'b000101, 6'b111111, 6'b111010, 6'b111000};
      end
   139: begin
        dout = {6'b001100, 6'b001000, 6'b111010, 6'b111001, 6'b111001, 6'b000100, 6'b001011, 6'b111101, 6'b110101, 6'b110111, 6'b111011, 6'b111001, 6'b000111, 6'b110001, 6'b110111, 6'b000100, 6'b000101, 6'b111100, 6'b110110, 6'b000101, 6'b110101, 6'b000110, 6'b000101, 6'b000110, 6'b111000, 6'b110101, 6'b110111, 6'b000101, 6'b000101, 6'b000101, 6'b000111, 6'b000110};
      end
   140: begin
        dout = {6'b111001, 6'b111000, 6'b000100, 6'b110110, 6'b110110, 6'b000011, 6'b110100, 6'b110101, 6'b110111, 6'b111000, 6'b110011, 6'b111000, 6'b110100, 6'b001000, 6'b110111, 6'b111111, 6'b110111, 6'b001011, 6'b001011, 6'b001001, 6'b111001, 6'b110010, 6'b110011, 6'b001011, 6'b110111, 6'b000101, 6'b110111, 6'b110100, 6'b111010, 6'b000011, 6'b111000, 6'b111010};
      end
   141: begin
        dout = {6'b001001, 6'b000110, 6'b000111, 6'b110100, 6'b000101, 6'b111011, 6'b001000, 6'b110010, 6'b000111, 6'b110000, 6'b001101, 6'b001001, 6'b110101, 6'b110011, 6'b001011, 6'b110110, 6'b111001, 6'b001010, 6'b000110, 6'b001010, 6'b000111, 6'b000011, 6'b111000, 6'b000111, 6'b000101, 6'b111100, 6'b110110, 6'b000110, 6'b110010, 6'b111100, 6'b110100, 6'b111101};
      end
   142: begin
        dout = {6'b001100, 6'b111011, 6'b110101, 6'b110111, 6'b001100, 6'b111011, 6'b001001, 6'b000110, 6'b110111, 6'b111000, 6'b000100, 6'b001001, 6'b110100, 6'b001101, 6'b000001, 6'b110100, 6'b000011, 6'b111010, 6'b110011, 6'b000100, 6'b110010, 6'b001101, 6'b001010, 6'b001101, 6'b111101, 6'b001000, 6'b000010, 6'b110111, 6'b000001, 6'b001010, 6'b101101, 6'b111001};
      end
   143: begin
        dout = {6'b001101, 6'b000010, 6'b000010, 6'b110110, 6'b111000, 6'b000101, 6'b000110, 6'b001100, 6'b001100, 6'b001110, 6'b110010, 6'b110111, 6'b001000, 6'b000011, 6'b110010, 6'b111010, 6'b000010, 6'b000101, 6'b000100, 6'b111010, 6'b110100, 6'b110000, 6'b110010, 6'b001000, 6'b111011, 6'b111100, 6'b000111, 6'b001001, 6'b001101, 6'b110100, 6'b111000, 6'b110110};
      end
   144: begin
        dout = {6'b001100, 6'b000100, 6'b000011, 6'b001000, 6'b001001, 6'b000011, 6'b000010, 6'b000110, 6'b111000, 6'b110111, 6'b001000, 6'b110101, 6'b001000, 6'b111100, 6'b000101, 6'b001110, 6'b110100, 6'b110111, 6'b001000, 6'b001101, 6'b000110, 6'b111001, 6'b000111, 6'b001100, 6'b000001, 6'b111100, 6'b000101, 6'b001011, 6'b110100, 6'b110111, 6'b111010, 6'b110110};
      end
   145: begin
        dout = {6'b110100, 6'b111011, 6'b000111, 6'b110010, 6'b000011, 6'b110110, 6'b000000, 6'b000001, 6'b000010, 6'b111110, 6'b001000, 6'b001000, 6'b111111, 6'b111110, 6'b000111, 6'b001010, 6'b001011, 6'b001000, 6'b001000, 6'b000011, 6'b001000, 6'b001001, 6'b001000, 6'b111101, 6'b110000, 6'b000101, 6'b000110, 6'b000101, 6'b110011, 6'b111110, 6'b001000, 6'b110111};
      end
   146: begin
        dout = {6'b110111, 6'b000111, 6'b000010, 6'b111011, 6'b001010, 6'b111001, 6'b000100, 6'b000100, 6'b111011, 6'b111010, 6'b000011, 6'b110110, 6'b111000, 6'b000101, 6'b110101, 6'b111000, 6'b000011, 6'b110101, 6'b000110, 6'b001100, 6'b000101, 6'b001100, 6'b000000, 6'b000011, 6'b111001, 6'b000101, 6'b000101, 6'b001001, 6'b000111, 6'b001101, 6'b001011, 6'b000010};
      end
   147: begin
        dout = {6'b111011, 6'b111011, 6'b001001, 6'b101101, 6'b110111, 6'b001110, 6'b000110, 6'b000111, 6'b001100, 6'b110100, 6'b001110, 6'b001101, 6'b111011, 6'b111000, 6'b000110, 6'b111100, 6'b001010, 6'b111001, 6'b111010, 6'b110011, 6'b001001, 6'b001010, 6'b111001, 6'b110100, 6'b111011, 6'b111011, 6'b000100, 6'b110111, 6'b001001, 6'b110110, 6'b001001, 6'b000101};
      end
   148: begin
        dout = {6'b001110, 6'b110110, 6'b001110, 6'b000101, 6'b000111, 6'b110110, 6'b111001, 6'b101111, 6'b001100, 6'b110111, 6'b110010, 6'b001011, 6'b000110, 6'b110110, 6'b001100, 6'b110000, 6'b001111, 6'b111011, 6'b110100, 6'b111111, 6'b110101, 6'b110111, 6'b111100, 6'b000101, 6'b000110, 6'b110110, 6'b000111, 6'b000111, 6'b001000, 6'b111010, 6'b110111, 6'b111000};
      end
   149: begin
        dout = {6'b110011, 6'b001000, 6'b111000, 6'b101111, 6'b111100, 6'b110101, 6'b111001, 6'b000011, 6'b111110, 6'b000100, 6'b000111, 6'b111010, 6'b110100, 6'b110011, 6'b001011, 6'b000110, 6'b111011, 6'b111011, 6'b111010, 6'b001011, 6'b001000, 6'b111011, 6'b110100, 6'b110110, 6'b110110, 6'b000000, 6'b111000, 6'b000000, 6'b111010, 6'b111111, 6'b000101, 6'b001000};
      end
   150: begin
        dout = {6'b110100, 6'b000101, 6'b111000, 6'b110010, 6'b110110, 6'b111000, 6'b111000, 6'b001110, 6'b111000, 6'b000110, 6'b000011, 6'b111100, 6'b111000, 6'b000100, 6'b111000, 6'b101111, 6'b001001, 6'b001001, 6'b110110, 6'b000101, 6'b110110, 6'b110110, 6'b111101, 6'b000011, 6'b110111, 6'b110110, 6'b110011, 6'b000110, 6'b110100, 6'b000011, 6'b001010, 6'b000011};
      end
   151: begin
        dout = {6'b110100, 6'b000101, 6'b110110, 6'b111010, 6'b111010, 6'b111101, 6'b110100, 6'b000011, 6'b110111, 6'b001110, 6'b111010, 6'b001111, 6'b111010, 6'b111100, 6'b111010, 6'b111010, 6'b110110, 6'b110100, 6'b001100, 6'b000111, 6'b111001, 6'b111011, 6'b111000, 6'b001010, 6'b001011, 6'b000110, 6'b001011, 6'b001000, 6'b001011, 6'b110111, 6'b111110, 6'b000111};
      end
   152: begin
        dout = {6'b000100, 6'b001000, 6'b000100, 6'b000111, 6'b000110, 6'b111000, 6'b110100, 6'b000110, 6'b000110, 6'b000001, 6'b000011, 6'b000010, 6'b110100, 6'b001010, 6'b000110, 6'b001001, 6'b110111, 6'b001101, 6'b000011, 6'b000110, 6'b110111, 6'b000101, 6'b111010, 6'b111110, 6'b000001, 6'b001000, 6'b000111, 6'b001000, 6'b110011, 6'b110101, 6'b101111, 6'b110111};
      end
   153: begin
        dout = {6'b001001, 6'b110010, 6'b000111, 6'b000111, 6'b111011, 6'b111000, 6'b110110, 6'b111010, 6'b001111, 6'b101110, 6'b010000, 6'b110110, 6'b001000, 6'b111001, 6'b000110, 6'b000101, 6'b110101, 6'b110111, 6'b000101, 6'b110101, 6'b001100, 6'b111011, 6'b001010, 6'b111001, 6'b111010, 6'b111010, 6'b000100, 6'b000000, 6'b110011, 6'b110111, 6'b111010, 6'b110100};
      end
   154: begin
        dout = {6'b110100, 6'b001001, 6'b000110, 6'b110101, 6'b000011, 6'b001000, 6'b000011, 6'b111110, 6'b000100, 6'b110011, 6'b110110, 6'b001010, 6'b110010, 6'b110101, 6'b110101, 6'b001000, 6'b110111, 6'b111000, 6'b110111, 6'b110110, 6'b111001, 6'b111010, 6'b110111, 6'b111110, 6'b110110, 6'b000001, 6'b110011, 6'b000111, 6'b001010, 6'b110111, 6'b110101, 6'b111010};
      end
   155: begin
        dout = {6'b110110, 6'b000111, 6'b000001, 6'b001111, 6'b000100, 6'b001000, 6'b001001, 6'b110111, 6'b000011, 6'b000111, 6'b001000, 6'b111010, 6'b111000, 6'b001011, 6'b111001, 6'b110101, 6'b110110, 6'b110000, 6'b000111, 6'b111101, 6'b000011, 6'b001000, 6'b010001, 6'b000110, 6'b111100, 6'b001010, 6'b000111, 6'b101110, 6'b110101, 6'b111101, 6'b110101, 6'b000101};
      end
   156: begin
        dout = {6'b110110, 6'b111011, 6'b110111, 6'b001010, 6'b110011, 6'b001100, 6'b110111, 6'b110111, 6'b111011, 6'b111001, 6'b000011, 6'b000110, 6'b110101, 6'b001000, 6'b111001, 6'b111011, 6'b110110, 6'b110100, 6'b000011, 6'b111011, 6'b110111, 6'b000110, 6'b001110, 6'b000110, 6'b110100, 6'b000100, 6'b001000, 6'b000110, 6'b001011, 6'b001001, 6'b001101, 6'b110000};
      end
   157: begin
        dout = {6'b110101, 6'b110100, 6'b001001, 6'b111010, 6'b000100, 6'b111110, 6'b110111, 6'b111010, 6'b000101, 6'b111110, 6'b001000, 6'b111000, 6'b111111, 6'b110010, 6'b000010, 6'b110100, 6'b000110, 6'b001100, 6'b001100, 6'b000111, 6'b001000, 6'b001011, 6'b001010, 6'b000011, 6'b000101, 6'b110100, 6'b001101, 6'b110110, 6'b001011, 6'b000101, 6'b111010, 6'b110111};
      end
   158: begin
        dout = {6'b111010, 6'b111100, 6'b001000, 6'b000001, 6'b000111, 6'b110010, 6'b001011, 6'b110011, 6'b111010, 6'b111010, 6'b001111, 6'b000110, 6'b001111, 6'b111001, 6'b001010, 6'b000111, 6'b001000, 6'b111000, 6'b001011, 6'b001100, 6'b110111, 6'b001000, 6'b001000, 6'b001001, 6'b001000, 6'b001000, 6'b001010, 6'b111011, 6'b001100, 6'b110010, 6'b000010, 6'b001000};
      end
   159: begin
        dout = {6'b111010, 6'b001101, 6'b111100, 6'b110101, 6'b000111, 6'b001000, 6'b111011, 6'b110111, 6'b111000, 6'b110100, 6'b000101, 6'b001001, 6'b111110, 6'b001101, 6'b110010, 6'b001010, 6'b110100, 6'b001001, 6'b000111, 6'b110111, 6'b111010, 6'b000101, 6'b001011, 6'b001110, 6'b111000, 6'b111011, 6'b000111, 6'b001001, 6'b111000, 6'b001000, 6'b000110, 6'b110111};
      end
   160: begin
        dout = {6'b111110, 6'b000100, 6'b000010, 6'b110011, 6'b000111, 6'b001011, 6'b110110, 6'b000100, 6'b001011, 6'b001011, 6'b000111, 6'b111010, 6'b110101, 6'b000111, 6'b000111, 6'b111001, 6'b110111, 6'b111110, 6'b000010, 6'b111000, 6'b110011, 6'b111001, 6'b000100, 6'b001011, 6'b000110, 6'b111010, 6'b001001, 6'b010000, 6'b000110, 6'b001110, 6'b000100, 6'b111001};
      end
   161: begin
        dout = {6'b111011, 6'b111010, 6'b001000, 6'b111010, 6'b000010, 6'b111001, 6'b111011, 6'b110011, 6'b000010, 6'b111001, 6'b110011, 6'b001000, 6'b000010, 6'b001101, 6'b111010, 6'b110001, 6'b000111, 6'b000110, 6'b001010, 6'b001000, 6'b001000, 6'b001100, 6'b111011, 6'b001000, 6'b110110, 6'b110110, 6'b000110, 6'b001001, 6'b111011, 6'b000101, 6'b000110, 6'b111011};
      end
   162: begin
        dout = {6'b111101, 6'b110101, 6'b110111, 6'b110111, 6'b000101, 6'b110100, 6'b111000, 6'b111000, 6'b111100, 6'b001001, 6'b111001, 6'b111001, 6'b110111, 6'b111001, 6'b110000, 6'b001111, 6'b001101, 6'b001010, 6'b000110, 6'b111010, 6'b000010, 6'b000100, 6'b000100, 6'b111010, 6'b111001, 6'b110110, 6'b110111, 6'b111100, 6'b001001, 6'b111001, 6'b110100, 6'b111010};
      end
   163: begin
        dout = {6'b111100, 6'b111100, 6'b101110, 6'b000101, 6'b000010, 6'b111000, 6'b001010, 6'b111101, 6'b110101, 6'b111110, 6'b110101, 6'b111000, 6'b111001, 6'b110101, 6'b001111, 6'b001010, 6'b001001, 6'b110111, 6'b111001, 6'b111000, 6'b000100, 6'b010010, 6'b110110, 6'b110110, 6'b110110, 6'b111000, 6'b000111, 6'b111011, 6'b111101, 6'b000101, 6'b101110, 6'b000111};
      end
   164: begin
        dout = {6'b110001, 6'b111001, 6'b000011, 6'b000111, 6'b010011, 6'b000100, 6'b110011, 6'b111101, 6'b000111, 6'b010001, 6'b111101, 6'b111100, 6'b110101, 6'b110110, 6'b111000, 6'b111001, 6'b111011, 6'b000010, 6'b000101, 6'b110101, 6'b001101, 6'b000100, 6'b111100, 6'b000111, 6'b000001, 6'b110000, 6'b001011, 6'b001001, 6'b000101, 6'b111001, 6'b110100, 6'b101110};
      end
   165: begin
        dout = {6'b111010, 6'b110100, 6'b110111, 6'b111111, 6'b111000, 6'b110100, 6'b000100, 6'b111101, 6'b001001, 6'b001110, 6'b110111, 6'b110101, 6'b000101, 6'b111001, 6'b001100, 6'b000111, 6'b000001, 6'b001101, 6'b111101, 6'b111100, 6'b000101, 6'b111100, 6'b111001, 6'b110110, 6'b110001, 6'b000100, 6'b111011, 6'b001001, 6'b000101, 6'b111001, 6'b001010, 6'b111000};
      end
   166: begin
        dout = {6'b001000, 6'b001001, 6'b000011, 6'b111001, 6'b111011, 6'b001100, 6'b000111, 6'b000001, 6'b110110, 6'b000101, 6'b111110, 6'b000100, 6'b111001, 6'b000100, 6'b111011, 6'b000001, 6'b000110, 6'b001001, 6'b111000, 6'b110100, 6'b111011, 6'b001010, 6'b001000, 6'b111100, 6'b001111, 6'b110100, 6'b000001, 6'b001110, 6'b111000, 6'b001100, 6'b110110, 6'b110111};
      end
   167: begin
        dout = {6'b110111, 6'b001100, 6'b000101, 6'b110110, 6'b000111, 6'b000110, 6'b000110, 6'b000111, 6'b001010, 6'b111100, 6'b110011, 6'b111000, 6'b110111, 6'b000111, 6'b000110, 6'b001101, 6'b110111, 6'b111001, 6'b111101, 6'b000001, 6'b000101, 6'b000100, 6'b111000, 6'b000100, 6'b001010, 6'b000101, 6'b110101, 6'b111010, 6'b111010, 6'b000001, 6'b111000, 6'b000110};
      end
   168: begin
        dout = {6'b111011, 6'b110111, 6'b000101, 6'b111011, 6'b001101, 6'b001000, 6'b001000, 6'b001000, 6'b111001, 6'b110001, 6'b111001, 6'b000101, 6'b110010, 6'b110110, 6'b111111, 6'b010001, 6'b000100, 6'b000110, 6'b111000, 6'b111100, 6'b111010, 6'b000110, 6'b110110, 6'b111000, 6'b111000, 6'b001000, 6'b000001, 6'b001000, 6'b001001, 6'b000111, 6'b111011, 6'b000110};
      end
   169: begin
        dout = {6'b000101, 6'b001010, 6'b110111, 6'b110110, 6'b110110, 6'b110110, 6'b001010, 6'b001000, 6'b111011, 6'b110101, 6'b110011, 6'b110111, 6'b111001, 6'b110110, 6'b001011, 6'b000000, 6'b001011, 6'b110111, 6'b001010, 6'b111000, 6'b000011, 6'b001011, 6'b110110, 6'b111100, 6'b110011, 6'b110010, 6'b110000, 6'b111010, 6'b001101, 6'b111001, 6'b110011, 6'b000111};
      end
   170: begin
        dout = {6'b001010, 6'b001000, 6'b001001, 6'b110110, 6'b110110, 6'b110110, 6'b110101, 6'b001000, 6'b111010, 6'b001001, 6'b000101, 6'b001111, 6'b110111, 6'b001000, 6'b000011, 6'b001010, 6'b000110, 6'b000100, 6'b000001, 6'b000101, 6'b000001, 6'b001001, 6'b111000, 6'b000011, 6'b111001, 6'b110111, 6'b001010, 6'b000111, 6'b000110, 6'b001001, 6'b000111, 6'b001000};
      end
   171: begin
        dout = {6'b111100, 6'b110111, 6'b001000, 6'b111000, 6'b001001, 6'b001000, 6'b111000, 6'b110111, 6'b110100, 6'b111001, 6'b110100, 6'b000101, 6'b110101, 6'b001100, 6'b110100, 6'b111001, 6'b111001, 6'b001001, 6'b110101, 6'b000010, 6'b110110, 6'b000110, 6'b001000, 6'b000101, 6'b001110, 6'b001101, 6'b111001, 6'b001101, 6'b111010, 6'b110011, 6'b001010, 6'b000110};
      end
   172: begin
        dout = {6'b001011, 6'b001000, 6'b000010, 6'b000110, 6'b000010, 6'b000100, 6'b001010, 6'b001100, 6'b001001, 6'b010001, 6'b000110, 6'b111011, 6'b110011, 6'b111100, 6'b101111, 6'b000101, 6'b111000, 6'b110111, 6'b110101, 6'b110101, 6'b110111, 6'b000111, 6'b110101, 6'b001011, 6'b111001, 6'b110111, 6'b110110, 6'b110110, 6'b110111, 6'b001010, 6'b001011, 6'b000011};
      end
   173: begin
        dout = {6'b001101, 6'b110111, 6'b001010, 6'b000111, 6'b111100, 6'b110101, 6'b000100, 6'b000111, 6'b110101, 6'b111010, 6'b000110, 6'b110101, 6'b111110, 6'b000010, 6'b111001, 6'b000111, 6'b111001, 6'b111001, 6'b001011, 6'b111010, 6'b111101, 6'b000110, 6'b001110, 6'b000110, 6'b000101, 6'b111110, 6'b000111, 6'b111000, 6'b110111, 6'b001100, 6'b000101, 6'b110000};
      end
   174: begin
        dout = {6'b001000, 6'b111011, 6'b000100, 6'b001010, 6'b000101, 6'b111001, 6'b110001, 6'b000110, 6'b000111, 6'b010000, 6'b000110, 6'b110010, 6'b110101, 6'b000101, 6'b001100, 6'b000100, 6'b001011, 6'b000110, 6'b111001, 6'b001010, 6'b001100, 6'b111101, 6'b111111, 6'b110100, 6'b000000, 6'b110111, 6'b110010, 6'b111010, 6'b000000, 6'b111110, 6'b111001, 6'b001001};
      end
   175: begin
        dout = {6'b001010, 6'b111000, 6'b111011, 6'b000110, 6'b000001, 6'b111100, 6'b110100, 6'b110100, 6'b001001, 6'b000101, 6'b001100, 6'b111000, 6'b111010, 6'b110110, 6'b110000, 6'b111010, 6'b111010, 6'b001100, 6'b000110, 6'b110011, 6'b110010, 6'b110011, 6'b110101, 6'b001001, 6'b001000, 6'b001001, 6'b001001, 6'b001001, 6'b000110, 6'b000100, 6'b111000, 6'b000010};
      end
   176: begin
        dout = {6'b001010, 6'b111011, 6'b110100, 6'b000101, 6'b111101, 6'b000011, 6'b000110, 6'b001001, 6'b110001, 6'b001100, 6'b001100, 6'b110100, 6'b001000, 6'b000111, 6'b110001, 6'b110111, 6'b000100, 6'b001001, 6'b001000, 6'b000110, 6'b000101, 6'b110111, 6'b110101, 6'b001011, 6'b110010, 6'b111000, 6'b001100, 6'b000110, 6'b111000, 6'b111010, 6'b000011, 6'b001000};
      end
   177: begin
        dout = {6'b110101, 6'b111011, 6'b000110, 6'b111000, 6'b110111, 6'b111011, 6'b001010, 6'b111001, 6'b001010, 6'b110111, 6'b110100, 6'b000110, 6'b110101, 6'b010001, 6'b111001, 6'b111001, 6'b010000, 6'b111100, 6'b001100, 6'b110111, 6'b000100, 6'b000011, 6'b111000, 6'b001000, 6'b000010, 6'b001010, 6'b111000, 6'b000111, 6'b000110, 6'b110011, 6'b001100, 6'b001111};
      end
   178: begin
        dout = {6'b000000, 6'b001001, 6'b000110, 6'b111000, 6'b110100, 6'b000111, 6'b110101, 6'b111010, 6'b110111, 6'b000101, 6'b111011, 6'b110011, 6'b111100, 6'b001111, 6'b111001, 6'b001011, 6'b000101, 6'b001100, 6'b000100, 6'b000111, 6'b001001, 6'b111000, 6'b110111, 6'b110101, 6'b001011, 6'b110111, 6'b000111, 6'b111001, 6'b000111, 6'b001010, 6'b001010, 6'b001001};
      end
   179: begin
        dout = {6'b111000, 6'b000111, 6'b110111, 6'b001110, 6'b000111, 6'b000101, 6'b001010, 6'b001000, 6'b110010, 6'b001000, 6'b001001, 6'b001101, 6'b001011, 6'b110100, 6'b001100, 6'b000110, 6'b110111, 6'b001100, 6'b000111, 6'b111010, 6'b111111, 6'b111100, 6'b000100, 6'b001100, 6'b001001, 6'b001000, 6'b110111, 6'b110001, 6'b000101, 6'b111100, 6'b111011, 6'b000111};
      end
   180: begin
        dout = {6'b000100, 6'b110111, 6'b110100, 6'b001011, 6'b110101, 6'b001101, 6'b111110, 6'b111111, 6'b001110, 6'b111111, 6'b110100, 6'b110101, 6'b111001, 6'b000100, 6'b000111, 6'b000010, 6'b110111, 6'b111110, 6'b001110, 6'b001000, 6'b110000, 6'b001001, 6'b110101, 6'b001001, 6'b111100, 6'b110111, 6'b000101, 6'b001000, 6'b001001, 6'b001000, 6'b111001, 6'b111001};
      end
   181: begin
        dout = {6'b111100, 6'b111010, 6'b000011, 6'b111010, 6'b111000, 6'b000110, 6'b000110, 6'b000101, 6'b001101, 6'b001011, 6'b111000, 6'b000111, 6'b111000, 6'b110111, 6'b111100, 6'b001001, 6'b000010, 6'b000111, 6'b110100, 6'b111000, 6'b000101, 6'b000111, 6'b111111, 6'b001001, 6'b001001, 6'b111000, 6'b110000, 6'b000101, 6'b111000, 6'b000111, 6'b111001, 6'b111100};
      end
   182: begin
        dout = {6'b110110, 6'b001110, 6'b000110, 6'b110011, 6'b001011, 6'b001000, 6'b000000, 6'b111100, 6'b001100, 6'b111010, 6'b111011, 6'b111100, 6'b110100, 6'b000000, 6'b111111, 6'b000011, 6'b001010, 6'b001001, 6'b001001, 6'b000100, 6'b000110, 6'b110110, 6'b001100, 6'b111101, 6'b111000, 6'b111101, 6'b001001, 6'b111000, 6'b001011, 6'b001000, 6'b000110, 6'b000100};
      end
   183: begin
        dout = {6'b000101, 6'b001100, 6'b110100, 6'b001100, 6'b000110, 6'b110111, 6'b111101, 6'b110110, 6'b110001, 6'b001001, 6'b001010, 6'b001010, 6'b111000, 6'b000110, 6'b001010, 6'b111101, 6'b111010, 6'b000100, 6'b111000, 6'b001000, 6'b001000, 6'b001000, 6'b000110, 6'b111100, 6'b001001, 6'b111001, 6'b000111, 6'b111000, 6'b000001, 6'b110110, 6'b111100, 6'b001010};
      end
   184: begin
        dout = {6'b001100, 6'b110010, 6'b001000, 6'b001001, 6'b110111, 6'b001011, 6'b001001, 6'b000111, 6'b000010, 6'b111011, 6'b000111, 6'b000001, 6'b000011, 6'b110101, 6'b101100, 6'b001110, 6'b110101, 6'b000000, 6'b110110, 6'b110101, 6'b001001, 6'b000101, 6'b110110, 6'b000111, 6'b110111, 6'b000100, 6'b111001, 6'b111000, 6'b110111, 6'b110110, 6'b110111, 6'b001010};
      end
   185: begin
        dout = {6'b000101, 6'b110111, 6'b001011, 6'b000110, 6'b000101, 6'b110111, 6'b001110, 6'b001001, 6'b111010, 6'b110100, 6'b000101, 6'b110011, 6'b111010, 6'b111011, 6'b111110, 6'b110111, 6'b110110, 6'b000011, 6'b000111, 6'b001010, 6'b111010, 6'b000011, 6'b001010, 6'b001101, 6'b000111, 6'b001101, 6'b001010, 6'b110101, 6'b111000, 6'b000100, 6'b000000, 6'b001100};
      end
   186: begin
        dout = {6'b000010, 6'b000011, 6'b000101, 6'b111110, 6'b000111, 6'b001100, 6'b000100, 6'b001111, 6'b111100, 6'b111000, 6'b001010, 6'b110001, 6'b110010, 6'b111011, 6'b010010, 6'b110110, 6'b111011, 6'b001000, 6'b000111, 6'b000110, 6'b000110, 6'b111011, 6'b000101, 6'b001000, 6'b001100, 6'b111000, 6'b111010, 6'b111111, 6'b111010, 6'b000111, 6'b000110, 6'b110110};
      end
   187: begin
        dout = {6'b110101, 6'b110100, 6'b000101, 6'b001001, 6'b111011, 6'b110110, 6'b111100, 6'b001001, 6'b001000, 6'b111111, 6'b111010, 6'b111000, 6'b111011, 6'b110100, 6'b111110, 6'b000110, 6'b110001, 6'b110101, 6'b001001, 6'b111001, 6'b111001, 6'b000011, 6'b110001, 6'b000100, 6'b000011, 6'b110011, 6'b000100, 6'b111011, 6'b001010, 6'b000100, 6'b110010, 6'b111010};
      end
   188: begin
        dout = {6'b110101, 6'b110001, 6'b000101, 6'b001001, 6'b111101, 6'b110110, 6'b001000, 6'b110100, 6'b111001, 6'b111010, 6'b111000, 6'b110111, 6'b111010, 6'b111010, 6'b110100, 6'b000100, 6'b000101, 6'b111010, 6'b001010, 6'b001000, 6'b110011, 6'b001100, 6'b110101, 6'b000111, 6'b110110, 6'b111010, 6'b001011, 6'b001011, 6'b000101, 6'b111010, 6'b110011, 6'b001111};
      end
   189: begin
        dout = {6'b111111, 6'b111000, 6'b000011, 6'b110101, 6'b110111, 6'b111000, 6'b001011, 6'b000110, 6'b001011, 6'b111000, 6'b000111, 6'b001100, 6'b000011, 6'b110110, 6'b000111, 6'b000110, 6'b110101, 6'b111101, 6'b111000, 6'b110010, 6'b000101, 6'b001011, 6'b001110, 6'b110100, 6'b001000, 6'b000001, 6'b111001, 6'b110101, 6'b110101, 6'b110101, 6'b111100, 6'b111001};
      end
   190: begin
        dout = {6'b111100, 6'b001110, 6'b111010, 6'b000111, 6'b000110, 6'b111010, 6'b111001, 6'b110101, 6'b001001, 6'b110110, 6'b000011, 6'b000111, 6'b001001, 6'b110100, 6'b110111, 6'b001101, 6'b000111, 6'b110111, 6'b111001, 6'b000010, 6'b111010, 6'b000110, 6'b111011, 6'b001000, 6'b110011, 6'b101101, 6'b111010, 6'b000000, 6'b000000, 6'b110101, 6'b000111, 6'b111100};
      end
   191: begin
        dout = {6'b001011, 6'b000011, 6'b000011, 6'b110000, 6'b110010, 6'b001100, 6'b001011, 6'b001010, 6'b110100, 6'b000100, 6'b110111, 6'b000011, 6'b111000, 6'b001010, 6'b001010, 6'b110111, 6'b111000, 6'b001011, 6'b110110, 6'b000011, 6'b111000, 6'b111010, 6'b110010, 6'b110011, 6'b000101, 6'b001010, 6'b000110, 6'b110101, 6'b001010, 6'b110010, 6'b001000, 6'b111011};
      end
   192: begin
        dout = {6'b000111, 6'b110101, 6'b111000, 6'b000110, 6'b000110, 6'b000011, 6'b110011, 6'b001001, 6'b000101, 6'b111111, 6'b110011, 6'b111011, 6'b111010, 6'b111010, 6'b110111, 6'b110011, 6'b110111, 6'b111010, 6'b000011, 6'b001010, 6'b001111, 6'b001011, 6'b110011, 6'b110101, 6'b110101, 6'b000011, 6'b000101, 6'b111010, 6'b111000, 6'b000100, 6'b000111, 6'b000101};
      end
   193: begin
        dout = {6'b001010, 6'b111000, 6'b111000, 6'b111000, 6'b110110, 6'b101111, 6'b001001, 6'b001010, 6'b001000, 6'b001011, 6'b001010, 6'b110100, 6'b000111, 6'b110101, 6'b111011, 6'b000101, 6'b001010, 6'b111100, 6'b111101, 6'b000101, 6'b110101, 6'b001100, 6'b001000, 6'b111011, 6'b000110, 6'b001011, 6'b111011, 6'b000111, 6'b001000, 6'b110100, 6'b000101, 6'b111001};
      end
   194: begin
        dout = {6'b111001, 6'b000011, 6'b001010, 6'b110111, 6'b000111, 6'b110011, 6'b000110, 6'b111100, 6'b001001, 6'b111010, 6'b110101, 6'b000111, 6'b111101, 6'b110010, 6'b000111, 6'b001000, 6'b110011, 6'b110110, 6'b111001, 6'b111011, 6'b110100, 6'b000111, 6'b000111, 6'b000010, 6'b111101, 6'b110100, 6'b000011, 6'b110100, 6'b110111, 6'b000111, 6'b111011, 6'b110110};
      end
   195: begin
        dout = {6'b000001, 6'b000010, 6'b110110, 6'b001010, 6'b111000, 6'b001011, 6'b001001, 6'b111010, 6'b111100, 6'b001100, 6'b001011, 6'b111100, 6'b000110, 6'b001100, 6'b110101, 6'b001100, 6'b111000, 6'b111100, 6'b111001, 6'b110110, 6'b000101, 6'b111000, 6'b111011, 6'b001000, 6'b110010, 6'b001010, 6'b000010, 6'b001101, 6'b111000, 6'b111110, 6'b110100, 6'b111111};
      end
   196: begin
        dout = {6'b000001, 6'b111011, 6'b000111, 6'b001000, 6'b111100, 6'b000100, 6'b000111, 6'b111000, 6'b110110, 6'b110101, 6'b000011, 6'b001001, 6'b110110, 6'b010000, 6'b111000, 6'b000110, 6'b111101, 6'b111100, 6'b000100, 6'b000011, 6'b001000, 6'b000110, 6'b111001, 6'b001000, 6'b110111, 6'b001101, 6'b111001, 6'b111110, 6'b001001, 6'b000101, 6'b110101, 6'b001000};
      end
   197: begin
        dout = {6'b001000, 6'b111010, 6'b111101, 6'b110100, 6'b111000, 6'b000111, 6'b110000, 6'b110110, 6'b001000, 6'b001000, 6'b001101, 6'b001011, 6'b001010, 6'b000101, 6'b111000, 6'b001000, 6'b110110, 6'b111011, 6'b110111, 6'b001011, 6'b000100, 6'b000001, 6'b001111, 6'b111001, 6'b110011, 6'b110100, 6'b111011, 6'b000101, 6'b001100, 6'b000110, 6'b000101, 6'b111001};
      end
   198: begin
        dout = {6'b001100, 6'b000101, 6'b000110, 6'b000100, 6'b110111, 6'b111011, 6'b000101, 6'b001101, 6'b000111, 6'b111101, 6'b111000, 6'b000101, 6'b110110, 6'b111011, 6'b110011, 6'b000100, 6'b001100, 6'b111111, 6'b000010, 6'b001100, 6'b001110, 6'b110111, 6'b001001, 6'b110011, 6'b111101, 6'b110101, 6'b110101, 6'b001100, 6'b000100, 6'b110101, 6'b111001, 6'b000101};
      end
   199: begin
        dout = {6'b000011, 6'b000011, 6'b110101, 6'b110101, 6'b000110, 6'b110100, 6'b111101, 6'b111101, 6'b110001, 6'b001011, 6'b110110, 6'b110110, 6'b000101, 6'b000100, 6'b111011, 6'b000110, 6'b001000, 6'b110011, 6'b001000, 6'b000011, 6'b000010, 6'b000010, 6'b110110, 6'b110011, 6'b001000, 6'b111100, 6'b000100, 6'b111010, 6'b001100, 6'b110011, 6'b001100, 6'b001100};
      end
   200: begin
        dout = {6'b111010, 6'b110111, 6'b000111, 6'b001101, 6'b000010, 6'b000110, 6'b110010, 6'b001101, 6'b110110, 6'b001001, 6'b000111, 6'b000101, 6'b111011, 6'b111001, 6'b110011, 6'b111000, 6'b000011, 6'b111001, 6'b001010, 6'b000100, 6'b001011, 6'b110110, 6'b000101, 6'b001000, 6'b001100, 6'b000110, 6'b101111, 6'b001100, 6'b001100, 6'b000011, 6'b001101, 6'b000100};
      end
   201: begin
        dout = {6'b000111, 6'b001000, 6'b111110, 6'b000001, 6'b110011, 6'b111011, 6'b000101, 6'b001001, 6'b000111, 6'b001010, 6'b110101, 6'b001100, 6'b111001, 6'b001110, 6'b110110, 6'b111000, 6'b111011, 6'b000101, 6'b110101, 6'b111000, 6'b110110, 6'b001000, 6'b001000, 6'b000100, 6'b001010, 6'b111010, 6'b000101, 6'b110111, 6'b001011, 6'b110110, 6'b110111, 6'b001010};
      end
   202: begin
        dout = {6'b111111, 6'b110101, 6'b000011, 6'b110110, 6'b000111, 6'b110111, 6'b000111, 6'b001010, 6'b110111, 6'b111000, 6'b110110, 6'b000101, 6'b000001, 6'b000000, 6'b000100, 6'b110000, 6'b111000, 6'b000110, 6'b000111, 6'b111001, 6'b111011, 6'b000111, 6'b110100, 6'b000001, 6'b001010, 6'b110100, 6'b111010, 6'b000100, 6'b110111, 6'b110100, 6'b001110, 6'b101111};
      end
   203: begin
        dout = {6'b001000, 6'b001101, 6'b000110, 6'b111001, 6'b001000, 6'b111111, 6'b001100, 6'b001001, 6'b110110, 6'b110100, 6'b000101, 6'b101110, 6'b000000, 6'b000110, 6'b111111, 6'b000100, 6'b000011, 6'b000000, 6'b111010, 6'b001111, 6'b111110, 6'b000111, 6'b001011, 6'b110101, 6'b110101, 6'b001110, 6'b111010, 6'b000110, 6'b111011, 6'b110110, 6'b000101, 6'b001000};
      end
   204: begin
        dout = {6'b110111, 6'b001101, 6'b001001, 6'b000101, 6'b110110, 6'b001010, 6'b000111, 6'b110110, 6'b001001, 6'b000110, 6'b110011, 6'b111011, 6'b110101, 6'b110110, 6'b001011, 6'b111100, 6'b000100, 6'b001000, 6'b000110, 6'b111010, 6'b110110, 6'b111100, 6'b111000, 6'b001010, 6'b110111, 6'b111101, 6'b110100, 6'b001000, 6'b110010, 6'b111011, 6'b110111, 6'b001100};
      end
   205: begin
        dout = {6'b000101, 6'b000111, 6'b000100, 6'b110101, 6'b111101, 6'b000110, 6'b000100, 6'b000100, 6'b001101, 6'b110110, 6'b001000, 6'b001101, 6'b000010, 6'b110111, 6'b111110, 6'b111011, 6'b110010, 6'b110100, 6'b110100, 6'b110100, 6'b111000, 6'b110110, 6'b000010, 6'b110111, 6'b000101, 6'b000101, 6'b001000, 6'b111010, 6'b001010, 6'b000101, 6'b000011, 6'b111001};
      end
   206: begin
        dout = {6'b000100, 6'b111100, 6'b000110, 6'b111001, 6'b110011, 6'b111001, 6'b001010, 6'b000100, 6'b001001, 6'b001010, 6'b111100, 6'b000011, 6'b110111, 6'b001010, 6'b001011, 6'b110011, 6'b000101, 6'b111000, 6'b000011, 6'b000111, 6'b001001, 6'b110010, 6'b001110, 6'b001000, 6'b000110, 6'b000111, 6'b111010, 6'b000111, 6'b001011, 6'b111101, 6'b111000, 6'b110011};
      end
   207: begin
        dout = {6'b001010, 6'b110011, 6'b000010, 6'b000110, 6'b001110, 6'b000110, 6'b001100, 6'b111011, 6'b000111, 6'b001001, 6'b000100, 6'b110110, 6'b000010, 6'b111111, 6'b001001, 6'b111010, 6'b111000, 6'b111000, 6'b111110, 6'b000011, 6'b110110, 6'b110001, 6'b001000, 6'b001110, 6'b111010, 6'b001010, 6'b111001, 6'b000100, 6'b000101, 6'b000101, 6'b111100, 6'b000011};
      end
   208: begin
        dout = {6'b001000, 6'b000010, 6'b000111, 6'b000110, 6'b110101, 6'b000011, 6'b001010, 6'b000111, 6'b001001, 6'b000100, 6'b000101, 6'b110011, 6'b110101, 6'b110010, 6'b111010, 6'b110111, 6'b111000, 6'b111010, 6'b001100, 6'b110111, 6'b001000, 6'b110011, 6'b000100, 6'b111011, 6'b110111, 6'b110010, 6'b000111, 6'b111011, 6'b111000, 6'b111010, 6'b001000, 6'b110101};
      end
   209: begin
        dout = {6'b010000, 6'b000110, 6'b111010, 6'b000000, 6'b110110, 6'b111000, 6'b001000, 6'b001010, 6'b110011, 6'b110110, 6'b111011, 6'b111000, 6'b111100, 6'b110101, 6'b110111, 6'b111001, 6'b110111, 6'b110110, 6'b111101, 6'b000111, 6'b111001, 6'b111011, 6'b111100, 6'b000101, 6'b000111, 6'b000100, 6'b110110, 6'b111100, 6'b111100, 6'b110101, 6'b110010, 6'b001011};
      end
   210: begin
        dout = {6'b110101, 6'b110110, 6'b110011, 6'b110100, 6'b001101, 6'b111000, 6'b111100, 6'b000111, 6'b000101, 6'b111110, 6'b001100, 6'b110110, 6'b110110, 6'b000011, 6'b000111, 6'b000111, 6'b000011, 6'b001010, 6'b110010, 6'b001001, 6'b001011, 6'b000001, 6'b001100, 6'b101110, 6'b110110, 6'b110011, 6'b110001, 6'b000100, 6'b110101, 6'b000000, 6'b001110, 6'b000100};
      end
   211: begin
        dout = {6'b110111, 6'b001000, 6'b000100, 6'b111000, 6'b001100, 6'b110110, 6'b001000, 6'b111100, 6'b111001, 6'b110001, 6'b001101, 6'b000101, 6'b110111, 6'b001010, 6'b001011, 6'b110100, 6'b111001, 6'b000110, 6'b110001, 6'b110110, 6'b110111, 6'b110101, 6'b001011, 6'b001111, 6'b111010, 6'b000001, 6'b001110, 6'b000110, 6'b110111, 6'b001000, 6'b110110, 6'b001011};
      end
   212: begin
        dout = {6'b001001, 6'b001001, 6'b111000, 6'b001001, 6'b000111, 6'b000111, 6'b001101, 6'b110110, 6'b110001, 6'b000010, 6'b001000, 6'b111100, 6'b111001, 6'b111010, 6'b111000, 6'b000100, 6'b111100, 6'b111000, 6'b111100, 6'b001000, 6'b111000, 6'b110111, 6'b000001, 6'b001011, 6'b001011, 6'b111000, 6'b110100, 6'b001101, 6'b111001, 6'b000010, 6'b111010, 6'b111011};
      end
   213: begin
        dout = {6'b111000, 6'b000111, 6'b001001, 6'b110011, 6'b110011, 6'b111011, 6'b001001, 6'b110110, 6'b111000, 6'b001000, 6'b111000, 6'b001110, 6'b110101, 6'b000110, 6'b000111, 6'b001100, 6'b110100, 6'b001011, 6'b001110, 6'b000000, 6'b111000, 6'b110110, 6'b001010, 6'b000101, 6'b111111, 6'b000011, 6'b110111, 6'b000111, 6'b001111, 6'b111011, 6'b000010, 6'b000000};
      end
   214: begin
        dout = {6'b001100, 6'b110110, 6'b111000, 6'b000011, 6'b110011, 6'b001111, 6'b001011, 6'b111000, 6'b000010, 6'b111011, 6'b001011, 6'b111000, 6'b000110, 6'b110100, 6'b111001, 6'b110011, 6'b000011, 6'b111000, 6'b001010, 6'b001010, 6'b000111, 6'b000111, 6'b000011, 6'b000110, 6'b001001, 6'b001000, 6'b110101, 6'b110100, 6'b000110, 6'b000001, 6'b000100, 6'b000011};
      end
   215: begin
        dout = {6'b000100, 6'b000110, 6'b111000, 6'b000111, 6'b111110, 6'b111010, 6'b110111, 6'b110011, 6'b000110, 6'b000011, 6'b111001, 6'b000001, 6'b110110, 6'b000101, 6'b000100, 6'b110110, 6'b001101, 6'b001010, 6'b000111, 6'b001001, 6'b000110, 6'b111011, 6'b111011, 6'b110100, 6'b111000, 6'b110001, 6'b110010, 6'b110110, 6'b001001, 6'b001001, 6'b111100, 6'b111001};
      end
   216: begin
        dout = {6'b111011, 6'b000001, 6'b001001, 6'b001001, 6'b001101, 6'b110100, 6'b111101, 6'b000100, 6'b110110, 6'b110011, 6'b110110, 6'b001100, 6'b001101, 6'b001001, 6'b001010, 6'b001010, 6'b110011, 6'b111010, 6'b110111, 6'b000101, 6'b001001, 6'b111000, 6'b111001, 6'b111010, 6'b110111, 6'b001001, 6'b111011, 6'b000101, 6'b000111, 6'b111001, 6'b111000, 6'b001111};
      end
   217: begin
        dout = {6'b110111, 6'b111000, 6'b111001, 6'b001111, 6'b001001, 6'b111001, 6'b111001, 6'b110101, 6'b001100, 6'b000101, 6'b111111, 6'b111001, 6'b111110, 6'b111110, 6'b111100, 6'b111011, 6'b111100, 6'b111001, 6'b000001, 6'b110110, 6'b001001, 6'b000101, 6'b110110, 6'b000111, 6'b110010, 6'b110001, 6'b001011, 6'b001010, 6'b110101, 6'b111001, 6'b000011, 6'b110001};
      end
   218: begin
        dout = {6'b110010, 6'b111010, 6'b111001, 6'b000101, 6'b110110, 6'b110101, 6'b110110, 6'b111001, 6'b000101, 6'b000111, 6'b000100, 6'b111111, 6'b111100, 6'b110110, 6'b001110, 6'b001010, 6'b000011, 6'b111000, 6'b000111, 6'b001011, 6'b000111, 6'b000010, 6'b110111, 6'b111010, 6'b001010, 6'b000100, 6'b000111, 6'b000010, 6'b000011, 6'b000110, 6'b001011, 6'b001011};
      end
   219: begin
        dout = {6'b111010, 6'b111001, 6'b001111, 6'b110110, 6'b000100, 6'b110111, 6'b110011, 6'b000100, 6'b110010, 6'b110110, 6'b000110, 6'b111011, 6'b111001, 6'b111000, 6'b001000, 6'b111011, 6'b110100, 6'b110101, 6'b001001, 6'b001001, 6'b111000, 6'b110000, 6'b110111, 6'b111011, 6'b000100, 6'b000100, 6'b110111, 6'b110010, 6'b110110, 6'b000110, 6'b000100, 6'b000111};
      end
   220: begin
        dout = {6'b001001, 6'b111001, 6'b110101, 6'b110110, 6'b110111, 6'b110000, 6'b111010, 6'b000110, 6'b111000, 6'b001010, 6'b001000, 6'b110111, 6'b110010, 6'b110100, 6'b111011, 6'b000000, 6'b110101, 6'b111011, 6'b001000, 6'b000011, 6'b110010, 6'b111101, 6'b001001, 6'b110101, 6'b000001, 6'b001010, 6'b000101, 6'b001000, 6'b111111, 6'b111001, 6'b001000, 6'b001000};
      end
   221: begin
        dout = {6'b000101, 6'b111011, 6'b101111, 6'b110100, 6'b001001, 6'b111101, 6'b111011, 6'b001011, 6'b001100, 6'b110011, 6'b110100, 6'b000101, 6'b000110, 6'b110101, 6'b001110, 6'b110100, 6'b111101, 6'b110111, 6'b001111, 6'b111101, 6'b111011, 6'b000101, 6'b001101, 6'b000110, 6'b001001, 6'b001000, 6'b111001, 6'b110111, 6'b110110, 6'b111000, 6'b110000, 6'b111010};
      end
   222: begin
        dout = {6'b111001, 6'b110100, 6'b000100, 6'b000111, 6'b001011, 6'b001011, 6'b110001, 6'b110111, 6'b110111, 6'b000010, 6'b001000, 6'b001100, 6'b111000, 6'b000101, 6'b111001, 6'b001011, 6'b001101, 6'b000101, 6'b111101, 6'b111001, 6'b000110, 6'b000011, 6'b110110, 6'b111000, 6'b000110, 6'b111100, 6'b111110, 6'b110110, 6'b111100, 6'b111110, 6'b000101, 6'b111100};
      end
   223: begin
        dout = {6'b001000, 6'b111000, 6'b001011, 6'b110000, 6'b111010, 6'b001001, 6'b111001, 6'b001010, 6'b101110, 6'b110111, 6'b111101, 6'b001001, 6'b111110, 6'b001011, 6'b111001, 6'b000110, 6'b000011, 6'b110110, 6'b001001, 6'b001000, 6'b111010, 6'b000110, 6'b000010, 6'b110111, 6'b000010, 6'b000110, 6'b000100, 6'b000011, 6'b000111, 6'b001010, 6'b110111, 6'b001111};
      end
   224: begin
        dout = {6'b000011, 6'b001000, 6'b001100, 6'b110100, 6'b110011, 6'b111001, 6'b110111, 6'b001110, 6'b110100, 6'b001010, 6'b001110, 6'b110100, 6'b000001, 6'b111000, 6'b001001, 6'b110110, 6'b001011, 6'b001101, 6'b110100, 6'b000101, 6'b001000, 6'b110101, 6'b001110, 6'b110111, 6'b110101, 6'b000111, 6'b111011, 6'b000110, 6'b000110, 6'b110101, 6'b110111, 6'b111000};
      end
   225: begin
        dout = {6'b000101, 6'b001000, 6'b111010, 6'b111011, 6'b000110, 6'b000110, 6'b111000, 6'b110111, 6'b110101, 6'b111010, 6'b110100, 6'b111010, 6'b110010, 6'b001011, 6'b001001, 6'b001001, 6'b000000, 6'b001011, 6'b110001, 6'b000100, 6'b110111, 6'b111010, 6'b000101, 6'b111000, 6'b010000, 6'b000000, 6'b110110, 6'b110011, 6'b000010, 6'b001110, 6'b111010, 6'b000011};
      end
   226: begin
        dout = {6'b111001, 6'b110101, 6'b111000, 6'b000001, 6'b111011, 6'b000001, 6'b111100, 6'b001010, 6'b001000, 6'b000111, 6'b111111, 6'b111101, 6'b000101, 6'b111001, 6'b111100, 6'b110101, 6'b111011, 6'b110101, 6'b111101, 6'b110100, 6'b110100, 6'b001010, 6'b001000, 6'b111101, 6'b110111, 6'b111110, 6'b001001, 6'b111000, 6'b111001, 6'b001100, 6'b000100, 6'b001001};
      end
   227: begin
        dout = {6'b110110, 6'b111011, 6'b110001, 6'b001000, 6'b000100, 6'b110010, 6'b110011, 6'b110101, 6'b111011, 6'b111000, 6'b001001, 6'b000100, 6'b001001, 6'b001101, 6'b001001, 6'b110110, 6'b111101, 6'b001100, 6'b110111, 6'b000100, 6'b111001, 6'b000010, 6'b001001, 6'b110100, 6'b111011, 6'b110101, 6'b001010, 6'b110110, 6'b001000, 6'b000111, 6'b001001, 6'b110111};
      end
   228: begin
        dout = {6'b000110, 6'b001000, 6'b001000, 6'b110110, 6'b001100, 6'b111010, 6'b110111, 6'b001001, 6'b000011, 6'b001000, 6'b111010, 6'b110110, 6'b010000, 6'b000111, 6'b110110, 6'b000010, 6'b111011, 6'b000111, 6'b001010, 6'b001000, 6'b110111, 6'b001010, 6'b001000, 6'b110100, 6'b110110, 6'b001011, 6'b000111, 6'b001011, 6'b000100, 6'b110100, 6'b111101, 6'b111011};
      end
   229: begin
        dout = {6'b110111, 6'b111110, 6'b111100, 6'b110110, 6'b111110, 6'b010010, 6'b110111, 6'b111010, 6'b111011, 6'b001011, 6'b000101, 6'b001001, 6'b000011, 6'b000001, 6'b110111, 6'b111000, 6'b000110, 6'b111010, 6'b000110, 6'b001011, 6'b001001, 6'b110001, 6'b110111, 6'b000111, 6'b111001, 6'b111101, 6'b111000, 6'b000111, 6'b001110, 6'b001100, 6'b001011, 6'b000110};
      end
   230: begin
        dout = {6'b001011, 6'b000100, 6'b001100, 6'b001111, 6'b110010, 6'b110111, 6'b110110, 6'b111000, 6'b110100, 6'b110111, 6'b000011, 6'b111000, 6'b000111, 6'b001000, 6'b001101, 6'b110110, 6'b000111, 6'b111011, 6'b000101, 6'b001100, 6'b111100, 6'b110101, 6'b111001, 6'b000011, 6'b110101, 6'b110110, 6'b110101, 6'b001100, 6'b000100, 6'b110111, 6'b111010, 6'b110101};
      end
   231: begin
        dout = {6'b001001, 6'b111011, 6'b110000, 6'b000100, 6'b000011, 6'b001001, 6'b001001, 6'b110010, 6'b110100, 6'b110111, 6'b111111, 6'b111001, 6'b111010, 6'b110101, 6'b000010, 6'b010000, 6'b110101, 6'b110100, 6'b111010, 6'b111011, 6'b000010, 6'b000111, 6'b000110, 6'b001010, 6'b000001, 6'b010010, 6'b111000, 6'b000100, 6'b110011, 6'b000011, 6'b110011, 6'b001101};
      end
   232: begin
        dout = {6'b001101, 6'b000011, 6'b000111, 6'b001000, 6'b111110, 6'b111100, 6'b110110, 6'b001110, 6'b000111, 6'b001100, 6'b001010, 6'b111100, 6'b000011, 6'b111101, 6'b001011, 6'b000011, 6'b000100, 6'b111001, 6'b110111, 6'b110011, 6'b111110, 6'b110110, 6'b000011, 6'b110100, 6'b111101, 6'b000000, 6'b001001, 6'b111000, 6'b001001, 6'b001111, 6'b000110, 6'b110100};
      end
   233: begin
        dout = {6'b110111, 6'b110100, 6'b111100, 6'b111100, 6'b001010, 6'b110011, 6'b001000, 6'b001001, 6'b001001, 6'b111101, 6'b001010, 6'b000101, 6'b110111, 6'b001110, 6'b110100, 6'b110100, 6'b111010, 6'b001100, 6'b001000, 6'b000111, 6'b111000, 6'b111001, 6'b001101, 6'b001000, 6'b001000, 6'b000110, 6'b110101, 6'b001011, 6'b000111, 6'b001000, 6'b000100, 6'b001000};
      end
   234: begin
        dout = {6'b111110, 6'b110100, 6'b001001, 6'b000000, 6'b001000, 6'b000100, 6'b111100, 6'b110101, 6'b000110, 6'b000101, 6'b111110, 6'b110100, 6'b111011, 6'b111010, 6'b001000, 6'b001010, 6'b111100, 6'b000111, 6'b110111, 6'b111010, 6'b110111, 6'b001100, 6'b001110, 6'b110111, 6'b000110, 6'b001000, 6'b000111, 6'b111101, 6'b001010, 6'b001010, 6'b000100, 6'b001100};
      end
   235: begin
        dout = {6'b001001, 6'b000001, 6'b001000, 6'b111010, 6'b001001, 6'b001100, 6'b111100, 6'b110100, 6'b110111, 6'b111101, 6'b110011, 6'b001000, 6'b111101, 6'b000100, 6'b000111, 6'b000001, 6'b000111, 6'b110100, 6'b110011, 6'b000110, 6'b000111, 6'b001001, 6'b000000, 6'b111011, 6'b001110, 6'b111010, 6'b111101, 6'b000011, 6'b110110, 6'b001110, 6'b000100, 6'b000110};
      end
   236: begin
        dout = {6'b000110, 6'b111010, 6'b001010, 6'b000111, 6'b110001, 6'b110010, 6'b001011, 6'b001011, 6'b000111, 6'b110111, 6'b110111, 6'b111101, 6'b000100, 6'b101111, 6'b110011, 6'b110110, 6'b110110, 6'b110011, 6'b111101, 6'b001010, 6'b110111, 6'b111010, 6'b001010, 6'b110111, 6'b111100, 6'b111101, 6'b000101, 6'b000111, 6'b111100, 6'b111101, 6'b110110, 6'b111011};
      end
   237: begin
        dout = {6'b000001, 6'b000110, 6'b000110, 6'b110010, 6'b110101, 6'b110101, 6'b010000, 6'b001010, 6'b000111, 6'b000000, 6'b000011, 6'b000100, 6'b000011, 6'b110011, 6'b001000, 6'b001000, 6'b110110, 6'b111100, 6'b111001, 6'b111011, 6'b010001, 6'b000101, 6'b110110, 6'b110110, 6'b001011, 6'b110000, 6'b101110, 6'b000100, 6'b110010, 6'b110101, 6'b110011, 6'b001001};
      end
   238: begin
        dout = {6'b001000, 6'b111000, 6'b110111, 6'b110110, 6'b001100, 6'b110011, 6'b000100, 6'b111100, 6'b001000, 6'b110101, 6'b000010, 6'b001011, 6'b110111, 6'b111010, 6'b110000, 6'b000001, 6'b000100, 6'b111101, 6'b110110, 6'b001000, 6'b111000, 6'b000010, 6'b001010, 6'b001111, 6'b001100, 6'b000011, 6'b110101, 6'b111101, 6'b001100, 6'b001010, 6'b000101, 6'b000000};
      end
   239: begin
        dout = {6'b110111, 6'b111001, 6'b000011, 6'b110101, 6'b111001, 6'b110111, 6'b000101, 6'b000100, 6'b110011, 6'b000111, 6'b111000, 6'b001010, 6'b111000, 6'b000110, 6'b111011, 6'b110101, 6'b110110, 6'b000111, 6'b000110, 6'b110111, 6'b111011, 6'b001000, 6'b001010, 6'b001100, 6'b001000, 6'b111011, 6'b000001, 6'b000111, 6'b111101, 6'b111010, 6'b111011, 6'b111011};
      end
   240: begin
        dout = {6'b111101, 6'b000110, 6'b111100, 6'b001001, 6'b111101, 6'b000111, 6'b110101, 6'b010000, 6'b001010, 6'b001001, 6'b001010, 6'b111000, 6'b000001, 6'b001110, 6'b110111, 6'b111001, 6'b000111, 6'b111100, 6'b000110, 6'b110000, 6'b001011, 6'b110010, 6'b001000, 6'b000111, 6'b001010, 6'b001000, 6'b001111, 6'b000011, 6'b001000, 6'b001001, 6'b001001, 6'b110110};
      end
   241: begin
        dout = {6'b110100, 6'b111100, 6'b000011, 6'b000100, 6'b000111, 6'b110111, 6'b001100, 6'b000101, 6'b000101, 6'b111011, 6'b111010, 6'b110100, 6'b000100, 6'b001010, 6'b111001, 6'b001011, 6'b000111, 6'b110010, 6'b000101, 6'b001000, 6'b001101, 6'b110010, 6'b110101, 6'b000111, 6'b001000, 6'b000101, 6'b000100, 6'b111001, 6'b110111, 6'b110010, 6'b001000, 6'b000001};
      end
   242: begin
        dout = {6'b001000, 6'b000110, 6'b001010, 6'b111011, 6'b000100, 6'b110011, 6'b111000, 6'b001010, 6'b110110, 6'b111010, 6'b000100, 6'b000101, 6'b111010, 6'b000111, 6'b110100, 6'b111010, 6'b001111, 6'b001011, 6'b111011, 6'b000111, 6'b110011, 6'b000110, 6'b111001, 6'b110101, 6'b111011, 6'b001110, 6'b000111, 6'b110100, 6'b001010, 6'b000111, 6'b111011, 6'b000100};
      end
   243: begin
        dout = {6'b110000, 6'b101111, 6'b000100, 6'b001000, 6'b111000, 6'b111011, 6'b001000, 6'b110101, 6'b000100, 6'b111001, 6'b000101, 6'b110111, 6'b000110, 6'b111011, 6'b111011, 6'b000101, 6'b000111, 6'b110100, 6'b000111, 6'b101101, 6'b111101, 6'b000101, 6'b110011, 6'b110011, 6'b111000, 6'b111001, 6'b111010, 6'b110111, 6'b110111, 6'b111000, 6'b000101, 6'b110101};
      end
   244: begin
        dout = {6'b111100, 6'b110101, 6'b000010, 6'b001001, 6'b001101, 6'b000001, 6'b001000, 6'b111110, 6'b000111, 6'b001110, 6'b001001, 6'b001101, 6'b001111, 6'b000001, 6'b111101, 6'b110110, 6'b001000, 6'b110110, 6'b111001, 6'b001010, 6'b111101, 6'b001001, 6'b110001, 6'b000010, 6'b111001, 6'b111011, 6'b000101, 6'b111010, 6'b110101, 6'b000110, 6'b001100, 6'b000100};
      end
   245: begin
        dout = {6'b110101, 6'b000110, 6'b110011, 6'b000000, 6'b010000, 6'b000100, 6'b001111, 6'b001101, 6'b110011, 6'b000111, 6'b110101, 6'b111101, 6'b111100, 6'b000111, 6'b111100, 6'b110101, 6'b110110, 6'b000000, 6'b111010, 6'b111000, 6'b000101, 6'b001000, 6'b110011, 6'b111110, 6'b001100, 6'b000001, 6'b111000, 6'b110111, 6'b001000, 6'b000101, 6'b111000, 6'b001100};
      end
   246: begin
        dout = {6'b111111, 6'b110100, 6'b000101, 6'b001001, 6'b000111, 6'b111011, 6'b000000, 6'b001100, 6'b001001, 6'b001110, 6'b000011, 6'b001001, 6'b110110, 6'b111010, 6'b110111, 6'b000101, 6'b110100, 6'b000010, 6'b110010, 6'b001100, 6'b001011, 6'b110100, 6'b000011, 6'b110101, 6'b111000, 6'b000100, 6'b110010, 6'b111010, 6'b110100, 6'b000110, 6'b111111, 6'b000111};
      end
   247: begin
        dout = {6'b001010, 6'b111100, 6'b000111, 6'b111001, 6'b001000, 6'b111101, 6'b111110, 6'b000101, 6'b110110, 6'b111011, 6'b110101, 6'b111001, 6'b000011, 6'b001000, 6'b111001, 6'b111011, 6'b001010, 6'b000100, 6'b000101, 6'b110101, 6'b000101, 6'b110100, 6'b000111, 6'b110001, 6'b001010, 6'b111000, 6'b001000, 6'b110111, 6'b001001, 6'b010000, 6'b111000, 6'b110110};
      end
   248: begin
        dout = {6'b111100, 6'b110001, 6'b110111, 6'b111000, 6'b110011, 6'b000100, 6'b000111, 6'b111001, 6'b111011, 6'b000000, 6'b111010, 6'b000011, 6'b111011, 6'b110011, 6'b001100, 6'b001110, 6'b001010, 6'b111000, 6'b110111, 6'b001100, 6'b001110, 6'b110110, 6'b001001, 6'b001000, 6'b000000, 6'b110001, 6'b001001, 6'b000010, 6'b111011, 6'b001010, 6'b110100, 6'b111010};
      end
   249: begin
        dout = {6'b111100, 6'b001000, 6'b111100, 6'b111001, 6'b101011, 6'b000111, 6'b000111, 6'b111010, 6'b000110, 6'b010000, 6'b110110, 6'b110110, 6'b111000, 6'b001100, 6'b111011, 6'b001001, 6'b110111, 6'b000010, 6'b111011, 6'b110100, 6'b110101, 6'b110101, 6'b111000, 6'b111101, 6'b111001, 6'b000101, 6'b000011, 6'b111110, 6'b110100, 6'b000101, 6'b111010, 6'b000110};
      end
   250: begin
        dout = {6'b000010, 6'b001000, 6'b110111, 6'b111100, 6'b000111, 6'b110000, 6'b110010, 6'b110101, 6'b001001, 6'b000011, 6'b001011, 6'b110110, 6'b110110, 6'b110110, 6'b000110, 6'b110100, 6'b110101, 6'b000101, 6'b001000, 6'b110101, 6'b110101, 6'b110110, 6'b111011, 6'b111000, 6'b000111, 6'b111011, 6'b110000, 6'b000110, 6'b111100, 6'b000000, 6'b110111, 6'b000101};
      end
   251: begin
        dout = {6'b001001, 6'b110110, 6'b111010, 6'b001011, 6'b111010, 6'b001000, 6'b000100, 6'b001101, 6'b110101, 6'b111010, 6'b110100, 6'b110100, 6'b001000, 6'b001011, 6'b110110, 6'b111000, 6'b000101, 6'b111001, 6'b110110, 6'b110110, 6'b001000, 6'b111001, 6'b111100, 6'b111110, 6'b000111, 6'b111000, 6'b001011, 6'b001110, 6'b001010, 6'b111000, 6'b001001, 6'b001101};
      end
   252: begin
        dout = {6'b000111, 6'b001001, 6'b000101, 6'b000101, 6'b111000, 6'b110001, 6'b111001, 6'b111001, 6'b110110, 6'b000110, 6'b110111, 6'b101101, 6'b111100, 6'b001100, 6'b000101, 6'b111001, 6'b111001, 6'b000100, 6'b111010, 6'b111000, 6'b110000, 6'b111101, 6'b111111, 6'b000010, 6'b110000, 6'b000111, 6'b110100, 6'b001001, 6'b110100, 6'b111011, 6'b111001, 6'b110100};
      end
   253: begin
        dout = {6'b111101, 6'b001101, 6'b000101, 6'b001100, 6'b111011, 6'b001010, 6'b001001, 6'b110001, 6'b000111, 6'b001001, 6'b001001, 6'b111011, 6'b001010, 6'b111001, 6'b110011, 6'b111010, 6'b110101, 6'b000100, 6'b110110, 6'b111001, 6'b000101, 6'b111111, 6'b111001, 6'b000101, 6'b001010, 6'b110110, 6'b111000, 6'b000101, 6'b110101, 6'b001011, 6'b110101, 6'b110010};
      end
   254: begin
        dout = {6'b001000, 6'b111011, 6'b110111, 6'b111000, 6'b111000, 6'b110101, 6'b111000, 6'b110111, 6'b111101, 6'b000100, 6'b110000, 6'b000111, 6'b110110, 6'b111001, 6'b000111, 6'b110000, 6'b000110, 6'b111010, 6'b111001, 6'b111000, 6'b001001, 6'b111001, 6'b000100, 6'b001000, 6'b111101, 6'b110001, 6'b110000, 6'b111110, 6'b001000, 6'b110011, 6'b001000, 6'b001001};
      end
   255: begin
        dout = {6'b111011, 6'b111011, 6'b001000, 6'b000110, 6'b110100, 6'b000010, 6'b001000, 6'b110110, 6'b001010, 6'b111111, 6'b111001, 6'b111000, 6'b110101, 6'b000011, 6'b110001, 6'b001010, 6'b111101, 6'b110111, 6'b110011, 6'b110111, 6'b000111, 6'b001000, 6'b110101, 6'b001100, 6'b111010, 6'b001010, 6'b001000, 6'b001000, 6'b101011, 6'b001101, 6'b001101, 6'b001000};
      end
   256: begin
        dout = {6'b110110, 6'b000110, 6'b000101, 6'b110111, 6'b111011, 6'b110101, 6'b110110, 6'b000001, 6'b111001, 6'b110010, 6'b101110, 6'b111100, 6'b000000, 6'b111101, 6'b111000, 6'b000110, 6'b110110, 6'b001101, 6'b111000, 6'b001010, 6'b111000, 6'b001010, 6'b000111, 6'b111011, 6'b110100, 6'b110111, 6'b111000, 6'b110100, 6'b001010, 6'b001000, 6'b001001, 6'b001011};
      end
   default: begin
        dout = {DW{1'b0}};
      end
 endcase
end//always
endmodule
