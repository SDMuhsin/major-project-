`timescale 1ns / 1ps
module Dmem_circ0_scripted(
		 muxOut,
		 dMemIn,
		 wr_en,
		 reaccessAddress,
		 reaccess_lyr,
		 rd_en, clk, rst 
 );
parameter r = 52;
parameter c = 13;
parameter w = 6;
parameter ADDRESSWIDTH = 5;

parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 
output wire [r*w -1 : 0]muxOut;// r numbers of w bits
input [r*w-1:0]dMemIn;
input wr_en;
input [ADDRESSWIDTH-1:0]reaccessAddress;
input reaccess_lyr;
input rd_en;
input clk,rst;

wire [(ADDRESSWIDTH+1)-1:0]case_sel;//{layer,address}
wire [w-1:0]dMemInDummy[r-1:0];
reg [w-1:0]muxOutWire[r-1:0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<r;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutWire[k];
        assign dMemInDummy[k] = dMemIn[ (k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always @(posedge clk) begin
    if (rst) begin
         for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] = 0;
           end
        end
    end
    else begin
    if(wr_en) begin
        // Set (i,j)th value = (i,j-1)th value
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Load Inputs
        for(i = r-1; i > -1; i=i-1) begin
            fifoOut[i][0] <= dMemInDummy[i]; 
        end
    end
    else begin 
        // Set (i,j)th value = (i,j)th value
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <= fifoOut[i][j];
            end
        end
    end
    end
end

assign case_sel = rd_en ? {reaccess_lyr,reaccessAddress} : {1'd1,READDISABLEDCASE};

always@(*) begin
    case(case_sel)

		 {1'd0, 5'd0} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd1} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd2} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd3} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd4} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd5} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd6} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd7} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 32 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 33 ][ 4 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 34 ][ 4 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 35 ][ 4 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 36 ][ 4 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 37 ][ 4 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 38 ][ 4 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 39 ][ 4 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 40 ][ 4 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 41 ][ 4 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 42 ][ 4 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 43 ][ 4 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 44 ][ 4 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 45 ][ 4 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 46 ][ 4 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 47 ][ 4 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 48 ][ 4 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 49 ][ 4 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 50 ][ 4 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd8} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 32 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 33 ][ 4 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 34 ][ 4 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 35 ][ 4 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 36 ][ 4 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 37 ][ 4 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 38 ][ 4 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 39 ][ 4 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 40 ][ 4 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 41 ][ 4 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 42 ][ 4 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 43 ][ 4 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 44 ][ 4 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 45 ][ 4 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 46 ][ 4 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 47 ][ 4 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 48 ][ 4 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 49 ][ 4 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 50 ][ 4 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd9} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 32 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 33 ][ 4 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 34 ][ 4 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 35 ][ 4 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 36 ][ 4 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 37 ][ 4 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 38 ][ 4 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 39 ][ 4 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 40 ][ 4 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 41 ][ 4 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 42 ][ 4 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 43 ][ 4 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 44 ][ 4 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 45 ][ 4 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 46 ][ 4 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 47 ][ 4 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 48 ][ 4 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 49 ][ 4 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 50 ][ 4 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd10} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 32 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 33 ][ 4 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 34 ][ 4 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 35 ][ 4 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 36 ][ 4 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 37 ][ 4 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 38 ][ 4 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 39 ][ 4 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 40 ][ 4 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 41 ][ 4 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 42 ][ 4 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 43 ][ 4 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 44 ][ 4 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 45 ][ 4 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 46 ][ 4 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 47 ][ 4 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 48 ][ 4 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 49 ][ 4 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 50 ][ 4 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd11} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 32 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 33 ][ 4 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 34 ][ 4 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 35 ][ 4 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 36 ][ 4 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 37 ][ 4 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 38 ][ 4 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 39 ][ 4 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 40 ][ 4 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 41 ][ 4 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 42 ][ 4 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 43 ][ 4 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 44 ][ 4 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 45 ][ 4 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 46 ][ 4 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 47 ][ 4 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 48 ][ 4 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 49 ][ 4 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 50 ][ 4 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd12} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 32 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 33 ][ 4 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 34 ][ 4 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 35 ][ 4 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 36 ][ 4 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 37 ][ 4 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 38 ][ 4 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 39 ][ 4 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 40 ][ 4 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 41 ][ 4 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 42 ][ 4 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 43 ][ 4 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 44 ][ 4 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 45 ][ 4 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 46 ][ 4 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 47 ][ 4 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 48 ][ 4 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 49 ][ 4 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 50 ][ 4 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = fifoOut[ 0 ][ 9 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 1 ][ 9 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 2 ][ 9 ]; 
		 end
		 {1'd0, 5'd13} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 32 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 33 ][ 4 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 34 ][ 4 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 35 ][ 4 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 36 ][ 4 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 37 ][ 4 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 38 ][ 4 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 39 ][ 4 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 40 ][ 4 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 41 ][ 4 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 42 ][ 4 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 43 ][ 4 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 44 ][ 4 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 45 ][ 4 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 46 ][ 4 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 47 ][ 4 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 48 ][ 4 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 49 ][ 4 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 50 ][ 4 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 3 ][ 10 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 4 ][ 10 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 5 ][ 10 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 6 ][ 10 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 7 ][ 10 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 8 ][ 10 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 9 ][ 10 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 10 ][ 10 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 11 ][ 10 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 12 ][ 10 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 13 ][ 10 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 14 ][ 10 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 15 ][ 10 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 16 ][ 10 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 17 ][ 10 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 18 ][ 10 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 19 ][ 10 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 20 ][ 10 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 21 ][ 10 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 22 ][ 10 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 23 ][ 10 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 24 ][ 10 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 25 ][ 10 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 0 ][ 9 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 1 ][ 9 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 2 ][ 9 ]; 
		 end
		 {1'd0, 5'd14} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 32 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 33 ][ 4 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 34 ][ 4 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 35 ][ 4 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 36 ][ 4 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 37 ][ 4 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 38 ][ 4 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 39 ][ 4 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 40 ][ 4 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 41 ][ 4 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 42 ][ 4 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 43 ][ 4 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 44 ][ 4 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 45 ][ 4 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 46 ][ 4 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 47 ][ 4 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 48 ][ 4 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 49 ][ 4 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 50 ][ 4 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 3 ][ 10 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 4 ][ 10 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 5 ][ 10 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 6 ][ 10 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 7 ][ 10 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 8 ][ 10 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 9 ][ 10 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 10 ][ 10 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 11 ][ 10 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 12 ][ 10 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 13 ][ 10 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 14 ][ 10 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 15 ][ 10 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 16 ][ 10 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 17 ][ 10 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 18 ][ 10 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 19 ][ 10 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 20 ][ 10 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 21 ][ 10 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 22 ][ 10 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 23 ][ 10 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 24 ][ 10 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 25 ][ 10 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 0 ][ 9 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 1 ][ 9 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 2 ][ 9 ]; 
		 end
		 {1'd0, 5'd15} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 32 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 33 ][ 4 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 34 ][ 4 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 35 ][ 4 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 36 ][ 4 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 37 ][ 4 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 38 ][ 4 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 39 ][ 4 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 40 ][ 4 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 41 ][ 4 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 42 ][ 4 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 43 ][ 4 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 44 ][ 4 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 45 ][ 4 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 46 ][ 4 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 47 ][ 4 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 48 ][ 4 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 49 ][ 4 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 50 ][ 4 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 3 ][ 10 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 4 ][ 10 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 5 ][ 10 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 6 ][ 10 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 7 ][ 10 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 8 ][ 10 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 9 ][ 10 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 10 ][ 10 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 11 ][ 10 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 12 ][ 10 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 13 ][ 10 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 14 ][ 10 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 15 ][ 10 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 16 ][ 10 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 17 ][ 10 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 18 ][ 10 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 19 ][ 10 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 20 ][ 10 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 21 ][ 10 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 22 ][ 10 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 23 ][ 10 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 24 ][ 10 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 25 ][ 10 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 0 ][ 9 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 1 ][ 9 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 2 ][ 9 ]; 
		 end
		 {1'd0, 5'd16} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 32 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 33 ][ 4 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 34 ][ 4 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 35 ][ 4 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 36 ][ 4 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 37 ][ 4 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 38 ][ 4 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 39 ][ 4 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 40 ][ 4 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 41 ][ 4 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 42 ][ 4 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 43 ][ 4 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 44 ][ 4 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 45 ][ 4 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 46 ][ 4 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 47 ][ 4 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 48 ][ 4 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 49 ][ 4 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 50 ][ 4 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 3 ][ 10 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 4 ][ 10 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 5 ][ 10 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 6 ][ 10 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 7 ][ 10 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 8 ][ 10 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 9 ][ 10 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 10 ][ 10 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 11 ][ 10 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 12 ][ 10 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 13 ][ 10 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 14 ][ 10 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 15 ][ 10 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 16 ][ 10 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 17 ][ 10 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 18 ][ 10 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 19 ][ 10 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 20 ][ 10 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 21 ][ 10 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 22 ][ 10 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 23 ][ 10 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 24 ][ 10 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 25 ][ 10 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 0 ][ 9 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 1 ][ 9 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 2 ][ 9 ]; 
		 end
		 {1'd0, 5'd17} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 32 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 33 ][ 4 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 34 ][ 4 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 35 ][ 4 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 36 ][ 4 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 37 ][ 4 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 38 ][ 4 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 39 ][ 4 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 40 ][ 4 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 41 ][ 4 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 42 ][ 4 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 43 ][ 4 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 44 ][ 4 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 45 ][ 4 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 46 ][ 4 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 47 ][ 4 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 48 ][ 4 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 49 ][ 4 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 50 ][ 4 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 3 ][ 10 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 4 ][ 10 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 5 ][ 10 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 6 ][ 10 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 7 ][ 10 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 8 ][ 10 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 9 ][ 10 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 10 ][ 10 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 11 ][ 10 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 12 ][ 10 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 13 ][ 10 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 14 ][ 10 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 15 ][ 10 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 16 ][ 10 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 17 ][ 10 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 18 ][ 10 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 19 ][ 10 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 20 ][ 10 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 21 ][ 10 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 22 ][ 10 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 23 ][ 10 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 24 ][ 10 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 25 ][ 10 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 0 ][ 9 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 1 ][ 9 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 2 ][ 9 ]; 
		 end
		 {1'd0, 5'd18} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 32 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 33 ][ 4 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 34 ][ 4 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 35 ][ 4 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 36 ][ 4 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 37 ][ 4 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 38 ][ 4 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 39 ][ 4 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 40 ][ 4 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 41 ][ 4 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 42 ][ 4 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 43 ][ 4 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 44 ][ 4 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 45 ][ 4 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 46 ][ 4 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 47 ][ 4 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 48 ][ 4 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 49 ][ 4 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 50 ][ 4 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 51 ][ 4 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 26 ][ 3 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 27 ][ 3 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 28 ][ 3 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 29 ][ 3 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 30 ][ 3 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 31 ][ 3 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 3 ][ 10 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 4 ][ 10 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 5 ][ 10 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 6 ][ 10 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 7 ][ 10 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 8 ][ 10 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 9 ][ 10 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 10 ][ 10 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 11 ][ 10 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 12 ][ 10 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 13 ][ 10 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 14 ][ 10 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 15 ][ 10 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 16 ][ 10 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 17 ][ 10 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 18 ][ 10 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 19 ][ 10 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 20 ][ 10 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 21 ][ 10 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 22 ][ 10 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 23 ][ 10 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 24 ][ 10 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 25 ][ 10 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 0 ][ 9 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 1 ][ 9 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 2 ][ 9 ]; 
		 end
		 {1'd0, 5'd19} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 32 ][ 4 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 33 ][ 4 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 34 ][ 4 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 35 ][ 4 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 36 ][ 4 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 37 ][ 4 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 38 ][ 4 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 39 ][ 4 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 40 ][ 4 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 41 ][ 4 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 42 ][ 4 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 43 ][ 4 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 44 ][ 4 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 45 ][ 4 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 46 ][ 4 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 47 ][ 4 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 48 ][ 4 ]; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 3 ][ 10 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 4 ][ 10 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 5 ][ 10 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 6 ][ 10 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 7 ][ 10 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 8 ][ 10 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 9 ][ 10 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 10 ][ 10 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 11 ][ 10 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 12 ][ 10 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 13 ][ 10 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 14 ][ 10 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 15 ][ 10 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 16 ][ 10 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 17 ][ 10 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 18 ][ 10 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 19 ][ 10 ]; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd0} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd1} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd2} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd3} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd4} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd5} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 8 ][ 2 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 9 ][ 2 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 10 ][ 2 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 11 ][ 2 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 12 ][ 2 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 13 ][ 2 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 14 ][ 2 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 15 ][ 2 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 16 ][ 2 ]; 
		 end
		 {1'd1, 5'd6} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 22 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 23 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 24 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 25 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 8 ][ 2 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 9 ][ 2 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 10 ][ 2 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 11 ][ 2 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 12 ][ 2 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 13 ][ 2 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 14 ][ 2 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 15 ][ 2 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 16 ][ 2 ]; 
		 end
		 {1'd1, 5'd7} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 22 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 23 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 24 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 25 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 8 ][ 2 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 9 ][ 2 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 10 ][ 2 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 11 ][ 2 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 12 ][ 2 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 13 ][ 2 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 14 ][ 2 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 15 ][ 2 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 16 ][ 2 ]; 
		 end
		 {1'd1, 5'd8} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 22 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 23 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 24 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 25 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 8 ][ 2 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 9 ][ 2 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 10 ][ 2 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 11 ][ 2 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 12 ][ 2 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 13 ][ 2 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 14 ][ 2 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 15 ][ 2 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 16 ][ 2 ]; 
		 end
		 {1'd1, 5'd9} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 22 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 23 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 24 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 25 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 8 ][ 2 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 9 ][ 2 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 10 ][ 2 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 11 ][ 2 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 12 ][ 2 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 13 ][ 2 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 14 ][ 2 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 15 ][ 2 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 16 ][ 2 ]; 
		 end
		 {1'd1, 5'd10} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 22 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 23 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 24 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 25 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 8 ][ 2 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 9 ][ 2 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 10 ][ 2 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 11 ][ 2 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 12 ][ 2 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 13 ][ 2 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 14 ][ 2 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 15 ][ 2 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 16 ][ 2 ]; 
		 end
		 {1'd1, 5'd11} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 22 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 23 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 24 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 25 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 8 ][ 2 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 9 ][ 2 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 10 ][ 2 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 11 ][ 2 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 12 ][ 2 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 13 ][ 2 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 14 ][ 2 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 15 ][ 2 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 16 ][ 2 ]; 
		 end
		 {1'd1, 5'd12} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 22 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 23 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 24 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 25 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 8 ][ 2 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 9 ][ 2 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 10 ][ 2 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 11 ][ 2 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 12 ][ 2 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 13 ][ 2 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 14 ][ 2 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 15 ][ 2 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 16 ][ 2 ]; 
		 end
		 {1'd1, 5'd13} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 22 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 23 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 24 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 25 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 8 ][ 2 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 9 ][ 2 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 10 ][ 2 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 11 ][ 2 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 12 ][ 2 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 13 ][ 2 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 14 ][ 2 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 15 ][ 2 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 16 ][ 2 ]; 
		 end
		 {1'd1, 5'd14} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = fifoOut[ 26 ][ 11 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 27 ][ 11 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 28 ][ 11 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 29 ][ 11 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 30 ][ 11 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 31 ][ 11 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 32 ][ 11 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 33 ][ 11 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 34 ][ 11 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 35 ][ 11 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 36 ][ 11 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 37 ][ 11 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 38 ][ 11 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 39 ][ 11 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 40 ][ 11 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 41 ][ 11 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 42 ][ 11 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 43 ][ 11 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 22 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 23 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 24 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 25 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 8 ][ 2 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 9 ][ 2 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 10 ][ 2 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 11 ][ 2 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 12 ][ 2 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 13 ][ 2 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 14 ][ 2 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 15 ][ 2 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 16 ][ 2 ]; 
		 end
		 {1'd1, 5'd15} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 44 ][ 12 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 45 ][ 12 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 46 ][ 12 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 47 ][ 12 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 48 ][ 12 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 49 ][ 12 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 50 ][ 12 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 51 ][ 12 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 26 ][ 11 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 27 ][ 11 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 28 ][ 11 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 29 ][ 11 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 30 ][ 11 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 31 ][ 11 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 32 ][ 11 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 33 ][ 11 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 34 ][ 11 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 35 ][ 11 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 36 ][ 11 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 37 ][ 11 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 38 ][ 11 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 39 ][ 11 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 40 ][ 11 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 41 ][ 11 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 42 ][ 11 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 43 ][ 11 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 22 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 23 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 24 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 25 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 8 ][ 2 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 9 ][ 2 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 10 ][ 2 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 11 ][ 2 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 12 ][ 2 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 13 ][ 2 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 14 ][ 2 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 15 ][ 2 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 16 ][ 2 ]; 
		 end
		 {1'd1, 5'd16} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 44 ][ 12 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 45 ][ 12 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 46 ][ 12 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 47 ][ 12 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 48 ][ 12 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 49 ][ 12 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 50 ][ 12 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 51 ][ 12 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 26 ][ 11 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 27 ][ 11 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 28 ][ 11 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 29 ][ 11 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 30 ][ 11 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 31 ][ 11 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 32 ][ 11 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 33 ][ 11 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 34 ][ 11 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 35 ][ 11 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 36 ][ 11 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 37 ][ 11 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 38 ][ 11 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 39 ][ 11 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 40 ][ 11 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 41 ][ 11 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 42 ][ 11 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 43 ][ 11 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 22 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 23 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 24 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 25 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 8 ][ 2 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 9 ][ 2 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 10 ][ 2 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 11 ][ 2 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 12 ][ 2 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 13 ][ 2 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 14 ][ 2 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 15 ][ 2 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 16 ][ 2 ]; 
		 end
		 {1'd1, 5'd17} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 44 ][ 12 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 45 ][ 12 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 46 ][ 12 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 47 ][ 12 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 48 ][ 12 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 49 ][ 12 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 50 ][ 12 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 51 ][ 12 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 26 ][ 11 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 27 ][ 11 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 28 ][ 11 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 29 ][ 11 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 30 ][ 11 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 31 ][ 11 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 32 ][ 11 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 33 ][ 11 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 34 ][ 11 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 35 ][ 11 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 36 ][ 11 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 37 ][ 11 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 38 ][ 11 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 39 ][ 11 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 40 ][ 11 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 41 ][ 11 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 42 ][ 11 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 43 ][ 11 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 22 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 23 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 24 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 25 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 8 ][ 2 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 9 ][ 2 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 10 ][ 2 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 11 ][ 2 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 12 ][ 2 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 13 ][ 2 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 14 ][ 2 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 15 ][ 2 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 16 ][ 2 ]; 
		 end
		 {1'd1, 5'd18} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 44 ][ 12 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 45 ][ 12 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 46 ][ 12 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 47 ][ 12 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 48 ][ 12 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 49 ][ 12 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 50 ][ 12 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 51 ][ 12 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 26 ][ 11 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 27 ][ 11 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 28 ][ 11 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 29 ][ 11 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 30 ][ 11 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 31 ][ 11 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 32 ][ 11 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 33 ][ 11 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 34 ][ 11 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 35 ][ 11 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 36 ][ 11 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 37 ][ 11 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 38 ][ 11 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 39 ][ 11 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 40 ][ 11 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 41 ][ 11 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 42 ][ 11 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 43 ][ 11 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 22 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 23 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 24 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 25 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 8 ][ 2 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 9 ][ 2 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 10 ][ 2 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 11 ][ 2 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 12 ][ 2 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 13 ][ 2 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 14 ][ 2 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 15 ][ 2 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 16 ][ 2 ]; 
		 end
		 {1'd1, 5'd19} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 44 ][ 12 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 45 ][ 12 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 46 ][ 12 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 47 ][ 12 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 48 ][ 12 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 49 ][ 12 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 50 ][ 12 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 51 ][ 12 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 26 ][ 11 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 27 ][ 11 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 28 ][ 11 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 29 ][ 11 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 30 ][ 11 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 31 ][ 11 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 32 ][ 11 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 33 ][ 11 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 34 ][ 11 ]; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 22 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 23 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 24 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 25 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 0 ][ 2 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 1 ][ 2 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 2 ][ 2 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 3 ][ 2 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 4 ][ 2 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 5 ][ 2 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 6 ][ 2 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 7 ][ 2 ]; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
    default:begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
    end
    endcase
end
endmodule
