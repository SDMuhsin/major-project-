`timescale 1ns / 1ps
module LMem1To0_511_circ7_yesshift_nounload_scripted(
        muxOut,
        ly0In,
        wr_en,
        feedback_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 11;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

input feedback_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        if(feedback_en) begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= fifoOut[i][c-1];
         end
        end
        else begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= ly0InConnector[i];
         end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[15][7];
              muxOutConnector[1] = fifoOut[16][7];
              muxOutConnector[2] = fifoOut[17][7];
              muxOutConnector[3] = fifoOut[18][7];
              muxOutConnector[4] = fifoOut[19][7];
              muxOutConnector[5] = fifoOut[20][7];
              muxOutConnector[6] = fifoOut[21][7];
              muxOutConnector[7] = fifoOut[22][7];
              muxOutConnector[8] = fifoOut[23][7];
              muxOutConnector[9] = fifoOut[24][7];
              muxOutConnector[10] = fifoOut[25][7];
              muxOutConnector[11] = fifoOut[0][6];
              muxOutConnector[12] = fifoOut[1][6];
              muxOutConnector[13] = fifoOut[2][6];
              muxOutConnector[14] = fifoOut[3][6];
              muxOutConnector[15] = fifoOut[4][6];
              muxOutConnector[16] = fifoOut[5][6];
              muxOutConnector[17] = fifoOut[6][6];
              muxOutConnector[18] = fifoOut[7][6];
              muxOutConnector[19] = fifoOut[8][6];
              muxOutConnector[20] = fifoOut[9][6];
              muxOutConnector[21] = fifoOut[10][6];
              muxOutConnector[22] = fifoOut[11][6];
              muxOutConnector[23] = fifoOut[12][6];
              muxOutConnector[24] = fifoOut[13][6];
              muxOutConnector[25] = fifoOut[14][6];
              muxOutConnector[26] = fifoOut[35][3];
              muxOutConnector[27] = fifoOut[36][3];
              muxOutConnector[28] = fifoOut[37][3];
              muxOutConnector[29] = fifoOut[38][3];
              muxOutConnector[30] = fifoOut[39][3];
              muxOutConnector[31] = fifoOut[40][3];
              muxOutConnector[32] = fifoOut[41][3];
              muxOutConnector[33] = fifoOut[42][3];
              muxOutConnector[34] = fifoOut[43][3];
              muxOutConnector[35] = fifoOut[44][3];
              muxOutConnector[36] = fifoOut[45][3];
              muxOutConnector[37] = fifoOut[46][3];
              muxOutConnector[38] = fifoOut[47][3];
              muxOutConnector[39] = fifoOut[48][3];
              muxOutConnector[40] = fifoOut[49][3];
              muxOutConnector[41] = fifoOut[50][3];
              muxOutConnector[42] = fifoOut[51][3];
              muxOutConnector[43] = fifoOut[26][2];
              muxOutConnector[44] = fifoOut[27][2];
              muxOutConnector[45] = fifoOut[28][2];
              muxOutConnector[46] = fifoOut[29][2];
              muxOutConnector[47] = fifoOut[30][2];
              muxOutConnector[48] = fifoOut[31][2];
              muxOutConnector[49] = fifoOut[32][2];
              muxOutConnector[50] = fifoOut[33][2];
              muxOutConnector[51] = fifoOut[34][2];
       end
       1: begin
              muxOutConnector[0] = fifoOut[15][7];
              muxOutConnector[1] = fifoOut[16][7];
              muxOutConnector[2] = fifoOut[17][7];
              muxOutConnector[3] = fifoOut[18][7];
              muxOutConnector[4] = fifoOut[19][7];
              muxOutConnector[5] = fifoOut[20][7];
              muxOutConnector[6] = fifoOut[21][7];
              muxOutConnector[7] = fifoOut[22][7];
              muxOutConnector[8] = fifoOut[23][7];
              muxOutConnector[9] = fifoOut[24][7];
              muxOutConnector[10] = fifoOut[25][7];
              muxOutConnector[11] = fifoOut[0][6];
              muxOutConnector[12] = fifoOut[1][6];
              muxOutConnector[13] = fifoOut[2][6];
              muxOutConnector[14] = fifoOut[3][6];
              muxOutConnector[15] = fifoOut[4][6];
              muxOutConnector[16] = fifoOut[5][6];
              muxOutConnector[17] = fifoOut[6][6];
              muxOutConnector[18] = fifoOut[7][6];
              muxOutConnector[19] = fifoOut[8][6];
              muxOutConnector[20] = fifoOut[9][6];
              muxOutConnector[21] = fifoOut[10][6];
              muxOutConnector[22] = fifoOut[11][6];
              muxOutConnector[23] = fifoOut[12][6];
              muxOutConnector[24] = fifoOut[13][6];
              muxOutConnector[25] = fifoOut[14][6];
              muxOutConnector[26] = fifoOut[35][3];
              muxOutConnector[27] = fifoOut[36][3];
              muxOutConnector[28] = fifoOut[37][3];
              muxOutConnector[29] = fifoOut[38][3];
              muxOutConnector[30] = fifoOut[39][3];
              muxOutConnector[31] = fifoOut[40][3];
              muxOutConnector[32] = fifoOut[41][3];
              muxOutConnector[33] = fifoOut[42][3];
              muxOutConnector[34] = fifoOut[43][3];
              muxOutConnector[35] = fifoOut[44][3];
              muxOutConnector[36] = fifoOut[45][3];
              muxOutConnector[37] = fifoOut[46][3];
              muxOutConnector[38] = fifoOut[47][3];
              muxOutConnector[39] = fifoOut[48][3];
              muxOutConnector[40] = fifoOut[49][3];
              muxOutConnector[41] = fifoOut[50][3];
              muxOutConnector[42] = fifoOut[51][3];
              muxOutConnector[43] = fifoOut[26][2];
              muxOutConnector[44] = fifoOut[27][2];
              muxOutConnector[45] = fifoOut[28][2];
              muxOutConnector[46] = fifoOut[29][2];
              muxOutConnector[47] = fifoOut[30][2];
              muxOutConnector[48] = fifoOut[31][2];
              muxOutConnector[49] = fifoOut[32][2];
              muxOutConnector[50] = fifoOut[33][2];
              muxOutConnector[51] = fifoOut[34][2];
       end
       2: begin
              muxOutConnector[0] = fifoOut[15][7];
              muxOutConnector[1] = fifoOut[16][7];
              muxOutConnector[2] = fifoOut[17][7];
              muxOutConnector[3] = fifoOut[18][7];
              muxOutConnector[4] = fifoOut[19][7];
              muxOutConnector[5] = fifoOut[20][7];
              muxOutConnector[6] = fifoOut[21][7];
              muxOutConnector[7] = fifoOut[22][7];
              muxOutConnector[8] = fifoOut[23][7];
              muxOutConnector[9] = fifoOut[24][7];
              muxOutConnector[10] = fifoOut[25][7];
              muxOutConnector[11] = fifoOut[0][6];
              muxOutConnector[12] = fifoOut[1][6];
              muxOutConnector[13] = fifoOut[2][6];
              muxOutConnector[14] = fifoOut[3][6];
              muxOutConnector[15] = fifoOut[4][6];
              muxOutConnector[16] = fifoOut[5][6];
              muxOutConnector[17] = fifoOut[6][6];
              muxOutConnector[18] = fifoOut[7][6];
              muxOutConnector[19] = fifoOut[8][6];
              muxOutConnector[20] = fifoOut[9][6];
              muxOutConnector[21] = fifoOut[10][6];
              muxOutConnector[22] = fifoOut[11][6];
              muxOutConnector[23] = fifoOut[12][6];
              muxOutConnector[24] = fifoOut[13][6];
              muxOutConnector[25] = fifoOut[14][6];
              muxOutConnector[26] = fifoOut[35][3];
              muxOutConnector[27] = fifoOut[36][3];
              muxOutConnector[28] = fifoOut[37][3];
              muxOutConnector[29] = fifoOut[38][3];
              muxOutConnector[30] = fifoOut[39][3];
              muxOutConnector[31] = fifoOut[40][3];
              muxOutConnector[32] = fifoOut[41][3];
              muxOutConnector[33] = fifoOut[42][3];
              muxOutConnector[34] = fifoOut[43][3];
              muxOutConnector[35] = fifoOut[44][3];
              muxOutConnector[36] = fifoOut[45][3];
              muxOutConnector[37] = fifoOut[46][3];
              muxOutConnector[38] = fifoOut[47][3];
              muxOutConnector[39] = fifoOut[48][3];
              muxOutConnector[40] = fifoOut[49][3];
              muxOutConnector[41] = fifoOut[50][3];
              muxOutConnector[42] = fifoOut[51][3];
              muxOutConnector[43] = fifoOut[26][2];
              muxOutConnector[44] = fifoOut[27][2];
              muxOutConnector[45] = fifoOut[28][2];
              muxOutConnector[46] = fifoOut[29][2];
              muxOutConnector[47] = fifoOut[30][2];
              muxOutConnector[48] = fifoOut[31][2];
              muxOutConnector[49] = fifoOut[32][2];
              muxOutConnector[50] = fifoOut[33][2];
              muxOutConnector[51] = fifoOut[34][2];
       end
       3: begin
              muxOutConnector[0] = fifoOut[15][7];
              muxOutConnector[1] = fifoOut[16][7];
              muxOutConnector[2] = fifoOut[17][7];
              muxOutConnector[3] = fifoOut[18][7];
              muxOutConnector[4] = fifoOut[19][7];
              muxOutConnector[5] = fifoOut[20][7];
              muxOutConnector[6] = fifoOut[21][7];
              muxOutConnector[7] = fifoOut[22][7];
              muxOutConnector[8] = fifoOut[23][7];
              muxOutConnector[9] = fifoOut[24][7];
              muxOutConnector[10] = fifoOut[25][7];
              muxOutConnector[11] = fifoOut[0][6];
              muxOutConnector[12] = fifoOut[1][6];
              muxOutConnector[13] = fifoOut[2][6];
              muxOutConnector[14] = fifoOut[3][6];
              muxOutConnector[15] = fifoOut[4][6];
              muxOutConnector[16] = fifoOut[5][6];
              muxOutConnector[17] = fifoOut[6][6];
              muxOutConnector[18] = fifoOut[7][6];
              muxOutConnector[19] = fifoOut[8][6];
              muxOutConnector[20] = fifoOut[9][6];
              muxOutConnector[21] = fifoOut[10][6];
              muxOutConnector[22] = fifoOut[11][6];
              muxOutConnector[23] = fifoOut[12][6];
              muxOutConnector[24] = fifoOut[13][6];
              muxOutConnector[25] = fifoOut[14][6];
              muxOutConnector[26] = fifoOut[35][3];
              muxOutConnector[27] = fifoOut[36][3];
              muxOutConnector[28] = fifoOut[37][3];
              muxOutConnector[29] = fifoOut[38][3];
              muxOutConnector[30] = fifoOut[39][3];
              muxOutConnector[31] = fifoOut[40][3];
              muxOutConnector[32] = fifoOut[41][3];
              muxOutConnector[33] = fifoOut[42][3];
              muxOutConnector[34] = fifoOut[18][2];
              muxOutConnector[35] = fifoOut[19][2];
              muxOutConnector[36] = fifoOut[20][2];
              muxOutConnector[37] = fifoOut[21][2];
              muxOutConnector[38] = fifoOut[22][2];
              muxOutConnector[39] = fifoOut[23][2];
              muxOutConnector[40] = fifoOut[24][2];
              muxOutConnector[41] = fifoOut[25][2];
              muxOutConnector[42] = fifoOut[0][1];
              muxOutConnector[43] = fifoOut[1][1];
              muxOutConnector[44] = fifoOut[2][1];
              muxOutConnector[45] = fifoOut[3][1];
              muxOutConnector[46] = fifoOut[4][1];
              muxOutConnector[47] = fifoOut[5][1];
              muxOutConnector[48] = fifoOut[6][1];
              muxOutConnector[49] = fifoOut[7][1];
              muxOutConnector[50] = fifoOut[8][1];
              muxOutConnector[51] = fifoOut[9][1];
       end
       4: begin
              muxOutConnector[0] = fifoOut[15][7];
              muxOutConnector[1] = fifoOut[16][7];
              muxOutConnector[2] = fifoOut[17][7];
              muxOutConnector[3] = fifoOut[18][7];
              muxOutConnector[4] = fifoOut[19][7];
              muxOutConnector[5] = fifoOut[20][7];
              muxOutConnector[6] = fifoOut[21][7];
              muxOutConnector[7] = fifoOut[22][7];
              muxOutConnector[8] = fifoOut[23][7];
              muxOutConnector[9] = fifoOut[24][7];
              muxOutConnector[10] = fifoOut[25][7];
              muxOutConnector[11] = fifoOut[0][6];
              muxOutConnector[12] = fifoOut[1][6];
              muxOutConnector[13] = fifoOut[2][6];
              muxOutConnector[14] = fifoOut[3][6];
              muxOutConnector[15] = fifoOut[4][6];
              muxOutConnector[16] = fifoOut[5][6];
              muxOutConnector[17] = fifoOut[6][6];
              muxOutConnector[18] = fifoOut[7][6];
              muxOutConnector[19] = fifoOut[8][6];
              muxOutConnector[20] = fifoOut[9][6];
              muxOutConnector[21] = fifoOut[10][6];
              muxOutConnector[22] = fifoOut[11][6];
              muxOutConnector[23] = fifoOut[12][6];
              muxOutConnector[24] = fifoOut[13][6];
              muxOutConnector[25] = fifoOut[14][6];
              muxOutConnector[26] = fifoOut[10][2];
              muxOutConnector[27] = fifoOut[11][2];
              muxOutConnector[28] = fifoOut[12][2];
              muxOutConnector[29] = fifoOut[13][2];
              muxOutConnector[30] = fifoOut[14][2];
              muxOutConnector[31] = fifoOut[15][2];
              muxOutConnector[32] = fifoOut[16][2];
              muxOutConnector[33] = fifoOut[17][2];
              muxOutConnector[34] = fifoOut[18][2];
              muxOutConnector[35] = fifoOut[19][2];
              muxOutConnector[36] = fifoOut[20][2];
              muxOutConnector[37] = fifoOut[21][2];
              muxOutConnector[38] = fifoOut[22][2];
              muxOutConnector[39] = fifoOut[23][2];
              muxOutConnector[40] = fifoOut[24][2];
              muxOutConnector[41] = fifoOut[25][2];
              muxOutConnector[42] = fifoOut[0][1];
              muxOutConnector[43] = fifoOut[1][1];
              muxOutConnector[44] = fifoOut[2][1];
              muxOutConnector[45] = fifoOut[3][1];
              muxOutConnector[46] = fifoOut[4][1];
              muxOutConnector[47] = fifoOut[5][1];
              muxOutConnector[48] = fifoOut[6][1];
              muxOutConnector[49] = fifoOut[7][1];
              muxOutConnector[50] = fifoOut[8][1];
              muxOutConnector[51] = fifoOut[9][1];
       end
       5: begin
              muxOutConnector[0] = fifoOut[15][7];
              muxOutConnector[1] = fifoOut[16][7];
              muxOutConnector[2] = fifoOut[17][7];
              muxOutConnector[3] = fifoOut[18][7];
              muxOutConnector[4] = fifoOut[19][7];
              muxOutConnector[5] = fifoOut[20][7];
              muxOutConnector[6] = fifoOut[21][7];
              muxOutConnector[7] = fifoOut[22][7];
              muxOutConnector[8] = fifoOut[23][7];
              muxOutConnector[9] = fifoOut[24][7];
              muxOutConnector[10] = fifoOut[25][7];
              muxOutConnector[11] = fifoOut[0][6];
              muxOutConnector[12] = fifoOut[1][6];
              muxOutConnector[13] = fifoOut[2][6];
              muxOutConnector[14] = fifoOut[3][6];
              muxOutConnector[15] = fifoOut[4][6];
              muxOutConnector[16] = fifoOut[5][6];
              muxOutConnector[17] = fifoOut[6][6];
              muxOutConnector[18] = fifoOut[7][6];
              muxOutConnector[19] = fifoOut[8][6];
              muxOutConnector[20] = fifoOut[9][6];
              muxOutConnector[21] = fifoOut[10][6];
              muxOutConnector[22] = fifoOut[11][6];
              muxOutConnector[23] = fifoOut[12][6];
              muxOutConnector[24] = fifoOut[13][6];
              muxOutConnector[25] = fifoOut[14][6];
              muxOutConnector[26] = fifoOut[10][2];
              muxOutConnector[27] = fifoOut[11][2];
              muxOutConnector[28] = fifoOut[12][2];
              muxOutConnector[29] = fifoOut[13][2];
              muxOutConnector[30] = fifoOut[14][2];
              muxOutConnector[31] = fifoOut[15][2];
              muxOutConnector[32] = fifoOut[16][2];
              muxOutConnector[33] = fifoOut[17][2];
              muxOutConnector[34] = fifoOut[18][2];
              muxOutConnector[35] = fifoOut[19][2];
              muxOutConnector[36] = fifoOut[20][2];
              muxOutConnector[37] = fifoOut[21][2];
              muxOutConnector[38] = fifoOut[22][2];
              muxOutConnector[39] = fifoOut[23][2];
              muxOutConnector[40] = fifoOut[24][2];
              muxOutConnector[41] = fifoOut[25][2];
              muxOutConnector[42] = fifoOut[0][1];
              muxOutConnector[43] = fifoOut[1][1];
              muxOutConnector[44] = fifoOut[2][1];
              muxOutConnector[45] = fifoOut[3][1];
              muxOutConnector[46] = fifoOut[4][1];
              muxOutConnector[47] = fifoOut[5][1];
              muxOutConnector[48] = fifoOut[6][1];
              muxOutConnector[49] = fifoOut[7][1];
              muxOutConnector[50] = fifoOut[8][1];
              muxOutConnector[51] = fifoOut[9][1];
       end
       6: begin
              muxOutConnector[0] = fifoOut[15][7];
              muxOutConnector[1] = fifoOut[16][7];
              muxOutConnector[2] = fifoOut[17][7];
              muxOutConnector[3] = fifoOut[18][7];
              muxOutConnector[4] = fifoOut[19][7];
              muxOutConnector[5] = fifoOut[20][7];
              muxOutConnector[6] = fifoOut[21][7];
              muxOutConnector[7] = fifoOut[22][7];
              muxOutConnector[8] = fifoOut[23][7];
              muxOutConnector[9] = fifoOut[24][7];
              muxOutConnector[10] = fifoOut[25][7];
              muxOutConnector[11] = fifoOut[0][6];
              muxOutConnector[12] = fifoOut[1][6];
              muxOutConnector[13] = fifoOut[2][6];
              muxOutConnector[14] = fifoOut[3][6];
              muxOutConnector[15] = fifoOut[4][6];
              muxOutConnector[16] = fifoOut[5][6];
              muxOutConnector[17] = fifoOut[6][6];
              muxOutConnector[18] = fifoOut[7][6];
              muxOutConnector[19] = fifoOut[8][6];
              muxOutConnector[20] = fifoOut[9][6];
              muxOutConnector[21] = fifoOut[10][6];
              muxOutConnector[22] = fifoOut[11][6];
              muxOutConnector[23] = fifoOut[12][6];
              muxOutConnector[24] = fifoOut[13][6];
              muxOutConnector[25] = fifoOut[14][6];
              muxOutConnector[26] = fifoOut[10][2];
              muxOutConnector[27] = fifoOut[11][2];
              muxOutConnector[28] = fifoOut[12][2];
              muxOutConnector[29] = fifoOut[13][2];
              muxOutConnector[30] = fifoOut[14][2];
              muxOutConnector[31] = fifoOut[15][2];
              muxOutConnector[32] = fifoOut[16][2];
              muxOutConnector[33] = fifoOut[17][2];
              muxOutConnector[34] = fifoOut[18][2];
              muxOutConnector[35] = fifoOut[19][2];
              muxOutConnector[36] = fifoOut[20][2];
              muxOutConnector[37] = fifoOut[21][2];
              muxOutConnector[38] = fifoOut[22][2];
              muxOutConnector[39] = fifoOut[23][2];
              muxOutConnector[40] = fifoOut[24][2];
              muxOutConnector[41] = fifoOut[25][2];
              muxOutConnector[42] = fifoOut[0][1];
              muxOutConnector[43] = fifoOut[1][1];
              muxOutConnector[44] = fifoOut[2][1];
              muxOutConnector[45] = fifoOut[3][1];
              muxOutConnector[46] = fifoOut[4][1];
              muxOutConnector[47] = fifoOut[5][1];
              muxOutConnector[48] = fifoOut[6][1];
              muxOutConnector[49] = fifoOut[7][1];
              muxOutConnector[50] = fifoOut[8][1];
              muxOutConnector[51] = fifoOut[9][1];
       end
       7: begin
              muxOutConnector[0] = fifoOut[15][7];
              muxOutConnector[1] = fifoOut[16][7];
              muxOutConnector[2] = fifoOut[51][6];
              muxOutConnector[3] = fifoOut[26][5];
              muxOutConnector[4] = fifoOut[27][5];
              muxOutConnector[5] = fifoOut[28][5];
              muxOutConnector[6] = fifoOut[29][5];
              muxOutConnector[7] = fifoOut[30][5];
              muxOutConnector[8] = fifoOut[31][5];
              muxOutConnector[9] = fifoOut[32][5];
              muxOutConnector[10] = fifoOut[33][5];
              muxOutConnector[11] = fifoOut[34][5];
              muxOutConnector[12] = fifoOut[35][5];
              muxOutConnector[13] = fifoOut[36][5];
              muxOutConnector[14] = fifoOut[37][5];
              muxOutConnector[15] = fifoOut[38][5];
              muxOutConnector[16] = fifoOut[39][5];
              muxOutConnector[17] = fifoOut[40][5];
              muxOutConnector[18] = fifoOut[41][5];
              muxOutConnector[19] = fifoOut[42][5];
              muxOutConnector[20] = fifoOut[43][5];
              muxOutConnector[21] = fifoOut[44][5];
              muxOutConnector[22] = fifoOut[45][5];
              muxOutConnector[23] = fifoOut[46][5];
              muxOutConnector[24] = fifoOut[47][5];
              muxOutConnector[25] = fifoOut[48][5];
              muxOutConnector[26] = fifoOut[10][2];
              muxOutConnector[27] = fifoOut[11][2];
              muxOutConnector[28] = fifoOut[12][2];
              muxOutConnector[29] = fifoOut[13][2];
              muxOutConnector[30] = fifoOut[14][2];
              muxOutConnector[31] = fifoOut[15][2];
              muxOutConnector[32] = fifoOut[16][2];
              muxOutConnector[33] = fifoOut[17][2];
              muxOutConnector[34] = fifoOut[18][2];
              muxOutConnector[35] = fifoOut[19][2];
              muxOutConnector[36] = fifoOut[20][2];
              muxOutConnector[37] = fifoOut[21][2];
              muxOutConnector[38] = fifoOut[22][2];
              muxOutConnector[39] = fifoOut[23][2];
              muxOutConnector[40] = fifoOut[24][2];
              muxOutConnector[41] = fifoOut[25][2];
              muxOutConnector[42] = fifoOut[0][1];
              muxOutConnector[43] = fifoOut[1][1];
              muxOutConnector[44] = fifoOut[2][1];
              muxOutConnector[45] = fifoOut[3][1];
              muxOutConnector[46] = fifoOut[4][1];
              muxOutConnector[47] = fifoOut[5][1];
              muxOutConnector[48] = fifoOut[6][1];
              muxOutConnector[49] = fifoOut[7][1];
              muxOutConnector[50] = fifoOut[8][1];
              muxOutConnector[51] = fifoOut[9][1];
       end
       8: begin
              muxOutConnector[0] = fifoOut[49][6];
              muxOutConnector[1] = fifoOut[50][6];
              muxOutConnector[2] = fifoOut[51][6];
              muxOutConnector[3] = fifoOut[26][5];
              muxOutConnector[4] = fifoOut[27][5];
              muxOutConnector[5] = fifoOut[28][5];
              muxOutConnector[6] = fifoOut[29][5];
              muxOutConnector[7] = fifoOut[30][5];
              muxOutConnector[8] = fifoOut[31][5];
              muxOutConnector[9] = fifoOut[32][5];
              muxOutConnector[10] = fifoOut[33][5];
              muxOutConnector[11] = fifoOut[34][5];
              muxOutConnector[12] = fifoOut[35][5];
              muxOutConnector[13] = fifoOut[36][5];
              muxOutConnector[14] = fifoOut[37][5];
              muxOutConnector[15] = fifoOut[38][5];
              muxOutConnector[16] = fifoOut[39][5];
              muxOutConnector[17] = fifoOut[40][5];
              muxOutConnector[18] = fifoOut[41][5];
              muxOutConnector[19] = fifoOut[42][5];
              muxOutConnector[20] = fifoOut[43][5];
              muxOutConnector[21] = fifoOut[44][5];
              muxOutConnector[22] = fifoOut[45][5];
              muxOutConnector[23] = fifoOut[46][5];
              muxOutConnector[24] = fifoOut[47][5];
              muxOutConnector[25] = fifoOut[48][5];
              muxOutConnector[26] = fifoOut[10][2];
              muxOutConnector[27] = fifoOut[11][2];
              muxOutConnector[28] = fifoOut[12][2];
              muxOutConnector[29] = fifoOut[13][2];
              muxOutConnector[30] = fifoOut[14][2];
              muxOutConnector[31] = fifoOut[15][2];
              muxOutConnector[32] = fifoOut[16][2];
              muxOutConnector[33] = fifoOut[17][2];
              muxOutConnector[34] = fifoOut[18][2];
              muxOutConnector[35] = fifoOut[19][2];
              muxOutConnector[36] = fifoOut[20][2];
              muxOutConnector[37] = fifoOut[21][2];
              muxOutConnector[38] = fifoOut[22][2];
              muxOutConnector[39] = fifoOut[23][2];
              muxOutConnector[40] = fifoOut[24][2];
              muxOutConnector[41] = fifoOut[25][2];
              muxOutConnector[42] = fifoOut[0][1];
              muxOutConnector[43] = fifoOut[1][1];
              muxOutConnector[44] = fifoOut[2][1];
              muxOutConnector[45] = fifoOut[3][1];
              muxOutConnector[46] = fifoOut[4][1];
              muxOutConnector[47] = fifoOut[5][1];
              muxOutConnector[48] = fifoOut[6][1];
              muxOutConnector[49] = fifoOut[7][1];
              muxOutConnector[50] = fifoOut[8][1];
              muxOutConnector[51] = fifoOut[9][1];
       end
       9: begin
              muxOutConnector[0] = fifoOut[49][6];
              muxOutConnector[1] = fifoOut[50][6];
              muxOutConnector[2] = fifoOut[51][6];
              muxOutConnector[3] = fifoOut[26][5];
              muxOutConnector[4] = fifoOut[27][5];
              muxOutConnector[5] = fifoOut[28][5];
              muxOutConnector[6] = fifoOut[29][5];
              muxOutConnector[7] = fifoOut[30][5];
              muxOutConnector[8] = fifoOut[31][5];
              muxOutConnector[9] = fifoOut[32][5];
              muxOutConnector[10] = fifoOut[33][5];
              muxOutConnector[11] = fifoOut[34][5];
              muxOutConnector[12] = fifoOut[35][5];
              muxOutConnector[13] = fifoOut[36][5];
              muxOutConnector[14] = fifoOut[37][5];
              muxOutConnector[15] = fifoOut[38][5];
              muxOutConnector[16] = fifoOut[39][5];
              muxOutConnector[17] = fifoOut[40][5];
              muxOutConnector[18] = fifoOut[41][5];
              muxOutConnector[19] = fifoOut[42][5];
              muxOutConnector[20] = fifoOut[43][5];
              muxOutConnector[21] = fifoOut[44][5];
              muxOutConnector[22] = fifoOut[45][5];
              muxOutConnector[23] = fifoOut[46][5];
              muxOutConnector[24] = fifoOut[47][5];
              muxOutConnector[25] = fifoOut[48][5];
              muxOutConnector[26] = fifoOut[10][2];
              muxOutConnector[27] = fifoOut[11][2];
              muxOutConnector[28] = fifoOut[12][2];
              muxOutConnector[29] = fifoOut[13][2];
              muxOutConnector[30] = fifoOut[14][2];
              muxOutConnector[31] = fifoOut[15][2];
              muxOutConnector[32] = fifoOut[16][2];
              muxOutConnector[33] = fifoOut[17][2];
              muxOutConnector[34] = fifoOut[18][2];
              muxOutConnector[35] = fifoOut[19][2];
              muxOutConnector[36] = fifoOut[20][2];
              muxOutConnector[37] = fifoOut[21][2];
              muxOutConnector[38] = fifoOut[22][2];
              muxOutConnector[39] = fifoOut[23][2];
              muxOutConnector[40] = fifoOut[24][2];
              muxOutConnector[41] = fifoOut[25][2];
              muxOutConnector[42] = fifoOut[0][1];
              muxOutConnector[43] = fifoOut[1][1];
              muxOutConnector[44] = fifoOut[2][1];
              muxOutConnector[45] = fifoOut[3][1];
              muxOutConnector[46] = fifoOut[4][1];
              muxOutConnector[47] = fifoOut[5][1];
              muxOutConnector[48] = fifoOut[6][1];
              muxOutConnector[49] = fifoOut[7][1];
              muxOutConnector[50] = fifoOut[8][1];
              muxOutConnector[51] = fifoOut[9][1];
       end
       10: begin
              muxOutConnector[0] = fifoOut[49][6];
              muxOutConnector[1] = fifoOut[50][6];
              muxOutConnector[2] = fifoOut[51][6];
              muxOutConnector[3] = fifoOut[26][5];
              muxOutConnector[4] = fifoOut[27][5];
              muxOutConnector[5] = fifoOut[28][5];
              muxOutConnector[6] = fifoOut[29][5];
              muxOutConnector[7] = fifoOut[30][5];
              muxOutConnector[8] = fifoOut[31][5];
              muxOutConnector[9] = fifoOut[32][5];
              muxOutConnector[10] = fifoOut[33][5];
              muxOutConnector[11] = fifoOut[34][5];
              muxOutConnector[12] = fifoOut[35][5];
              muxOutConnector[13] = fifoOut[36][5];
              muxOutConnector[14] = fifoOut[37][5];
              muxOutConnector[15] = fifoOut[38][5];
              muxOutConnector[16] = fifoOut[39][5];
              muxOutConnector[17] = fifoOut[40][5];
              muxOutConnector[18] = fifoOut[41][5];
              muxOutConnector[19] = fifoOut[42][5];
              muxOutConnector[20] = fifoOut[43][5];
              muxOutConnector[21] = fifoOut[44][5];
              muxOutConnector[22] = fifoOut[45][5];
              muxOutConnector[23] = fifoOut[46][5];
              muxOutConnector[24] = fifoOut[47][5];
              muxOutConnector[25] = fifoOut[48][5];
              muxOutConnector[26] = fifoOut[10][2];
              muxOutConnector[27] = fifoOut[11][2];
              muxOutConnector[28] = fifoOut[12][2];
              muxOutConnector[29] = fifoOut[13][2];
              muxOutConnector[30] = fifoOut[14][2];
              muxOutConnector[31] = fifoOut[15][2];
              muxOutConnector[32] = fifoOut[16][2];
              muxOutConnector[33] = fifoOut[17][2];
              muxOutConnector[34] = fifoOut[18][2];
              muxOutConnector[35] = fifoOut[19][2];
              muxOutConnector[36] = fifoOut[20][2];
              muxOutConnector[37] = fifoOut[21][2];
              muxOutConnector[38] = fifoOut[22][2];
              muxOutConnector[39] = fifoOut[23][2];
              muxOutConnector[40] = fifoOut[24][2];
              muxOutConnector[41] = fifoOut[25][2];
              muxOutConnector[42] = fifoOut[0][1];
              muxOutConnector[43] = fifoOut[1][1];
              muxOutConnector[44] = fifoOut[2][1];
              muxOutConnector[45] = fifoOut[3][1];
              muxOutConnector[46] = fifoOut[4][1];
              muxOutConnector[47] = fifoOut[5][1];
              muxOutConnector[48] = fifoOut[6][1];
              muxOutConnector[49] = fifoOut[7][1];
              muxOutConnector[50] = fifoOut[8][1];
              muxOutConnector[51] = fifoOut[9][1];
       end
       11: begin
              muxOutConnector[0] = fifoOut[49][6];
              muxOutConnector[1] = fifoOut[50][6];
              muxOutConnector[2] = fifoOut[51][6];
              muxOutConnector[3] = fifoOut[26][5];
              muxOutConnector[4] = fifoOut[27][5];
              muxOutConnector[5] = fifoOut[28][5];
              muxOutConnector[6] = fifoOut[29][5];
              muxOutConnector[7] = fifoOut[30][5];
              muxOutConnector[8] = fifoOut[31][5];
              muxOutConnector[9] = fifoOut[32][5];
              muxOutConnector[10] = fifoOut[33][5];
              muxOutConnector[11] = fifoOut[34][5];
              muxOutConnector[12] = fifoOut[35][5];
              muxOutConnector[13] = fifoOut[36][5];
              muxOutConnector[14] = fifoOut[37][5];
              muxOutConnector[15] = fifoOut[38][5];
              muxOutConnector[16] = fifoOut[39][5];
              muxOutConnector[17] = fifoOut[40][5];
              muxOutConnector[18] = fifoOut[41][5];
              muxOutConnector[19] = fifoOut[42][5];
              muxOutConnector[20] = fifoOut[43][5];
              muxOutConnector[21] = fifoOut[44][5];
              muxOutConnector[22] = fifoOut[45][5];
              muxOutConnector[23] = fifoOut[46][5];
              muxOutConnector[24] = fifoOut[47][5];
              muxOutConnector[25] = fifoOut[48][5];
              muxOutConnector[26] = fifoOut[10][2];
              muxOutConnector[27] = fifoOut[11][2];
              muxOutConnector[28] = fifoOut[12][2];
              muxOutConnector[29] = fifoOut[13][2];
              muxOutConnector[30] = fifoOut[14][2];
              muxOutConnector[31] = fifoOut[15][2];
              muxOutConnector[32] = fifoOut[16][2];
              muxOutConnector[33] = fifoOut[17][2];
              muxOutConnector[34] = fifoOut[18][2];
              muxOutConnector[35] = fifoOut[19][2];
              muxOutConnector[36] = fifoOut[20][2];
              muxOutConnector[37] = fifoOut[21][2];
              muxOutConnector[38] = fifoOut[22][2];
              muxOutConnector[39] = fifoOut[23][2];
              muxOutConnector[40] = fifoOut[24][2];
              muxOutConnector[41] = fifoOut[25][2];
              muxOutConnector[42] = fifoOut[0][1];
              muxOutConnector[43] = fifoOut[1][1];
              muxOutConnector[44] = fifoOut[2][1];
              muxOutConnector[45] = fifoOut[3][1];
              muxOutConnector[46] = fifoOut[4][1];
              muxOutConnector[47] = fifoOut[5][1];
              muxOutConnector[48] = fifoOut[6][1];
              muxOutConnector[49] = fifoOut[7][1];
              muxOutConnector[50] = fifoOut[8][1];
              muxOutConnector[51] = fifoOut[9][1];
       end
       12: begin
              muxOutConnector[0] = fifoOut[49][6];
              muxOutConnector[1] = fifoOut[50][6];
              muxOutConnector[2] = fifoOut[51][6];
              muxOutConnector[3] = fifoOut[26][5];
              muxOutConnector[4] = fifoOut[27][5];
              muxOutConnector[5] = fifoOut[28][5];
              muxOutConnector[6] = fifoOut[29][5];
              muxOutConnector[7] = fifoOut[30][5];
              muxOutConnector[8] = fifoOut[31][5];
              muxOutConnector[9] = fifoOut[32][5];
              muxOutConnector[10] = fifoOut[33][5];
              muxOutConnector[11] = fifoOut[34][5];
              muxOutConnector[12] = fifoOut[35][5];
              muxOutConnector[13] = fifoOut[36][5];
              muxOutConnector[14] = fifoOut[37][5];
              muxOutConnector[15] = fifoOut[38][5];
              muxOutConnector[16] = fifoOut[39][5];
              muxOutConnector[17] = fifoOut[40][5];
              muxOutConnector[18] = fifoOut[41][5];
              muxOutConnector[19] = fifoOut[42][5];
              muxOutConnector[20] = fifoOut[43][5];
              muxOutConnector[21] = fifoOut[44][5];
              muxOutConnector[22] = fifoOut[45][5];
              muxOutConnector[23] = fifoOut[46][5];
              muxOutConnector[24] = fifoOut[47][5];
              muxOutConnector[25] = fifoOut[48][5];
              muxOutConnector[26] = fifoOut[10][2];
              muxOutConnector[27] = fifoOut[11][2];
              muxOutConnector[28] = fifoOut[12][2];
              muxOutConnector[29] = fifoOut[13][2];
              muxOutConnector[30] = fifoOut[14][2];
              muxOutConnector[31] = fifoOut[15][2];
              muxOutConnector[32] = fifoOut[16][2];
              muxOutConnector[33] = fifoOut[17][2];
              muxOutConnector[34] = fifoOut[18][2];
              muxOutConnector[35] = fifoOut[19][2];
              muxOutConnector[36] = fifoOut[20][2];
              muxOutConnector[37] = fifoOut[21][2];
              muxOutConnector[38] = fifoOut[22][2];
              muxOutConnector[39] = fifoOut[23][2];
              muxOutConnector[40] = fifoOut[24][2];
              muxOutConnector[41] = fifoOut[25][2];
              muxOutConnector[42] = fifoOut[0][1];
              muxOutConnector[43] = fifoOut[1][1];
              muxOutConnector[44] = fifoOut[2][1];
              muxOutConnector[45] = fifoOut[3][1];
              muxOutConnector[46] = fifoOut[4][1];
              muxOutConnector[47] = fifoOut[5][1];
              muxOutConnector[48] = fifoOut[6][1];
              muxOutConnector[49] = fifoOut[7][1];
              muxOutConnector[50] = fifoOut[8][1];
              muxOutConnector[51] = fifoOut[9][1];
       end
       13: begin
              muxOutConnector[0] = fifoOut[49][6];
              muxOutConnector[1] = fifoOut[50][6];
              muxOutConnector[2] = fifoOut[51][6];
              muxOutConnector[3] = fifoOut[26][5];
              muxOutConnector[4] = fifoOut[27][5];
              muxOutConnector[5] = fifoOut[28][5];
              muxOutConnector[6] = fifoOut[29][5];
              muxOutConnector[7] = fifoOut[30][5];
              muxOutConnector[8] = fifoOut[31][5];
              muxOutConnector[9] = fifoOut[32][5];
              muxOutConnector[10] = fifoOut[33][5];
              muxOutConnector[11] = fifoOut[34][5];
              muxOutConnector[12] = fifoOut[35][5];
              muxOutConnector[13] = fifoOut[36][5];
              muxOutConnector[14] = fifoOut[37][5];
              muxOutConnector[15] = fifoOut[38][5];
              muxOutConnector[16] = fifoOut[39][5];
              muxOutConnector[17] = fifoOut[40][5];
              muxOutConnector[18] = fifoOut[41][5];
              muxOutConnector[19] = fifoOut[42][5];
              muxOutConnector[20] = fifoOut[43][5];
              muxOutConnector[21] = fifoOut[44][5];
              muxOutConnector[22] = fifoOut[45][5];
              muxOutConnector[23] = fifoOut[46][5];
              muxOutConnector[24] = fifoOut[47][5];
              muxOutConnector[25] = fifoOut[48][5];
              muxOutConnector[26] = fifoOut[10][2];
              muxOutConnector[27] = fifoOut[11][2];
              muxOutConnector[28] = fifoOut[12][2];
              muxOutConnector[29] = fifoOut[13][2];
              muxOutConnector[30] = fifoOut[14][2];
              muxOutConnector[31] = fifoOut[15][2];
              muxOutConnector[32] = fifoOut[16][2];
              muxOutConnector[33] = fifoOut[51][1];
              muxOutConnector[34] = fifoOut[26][0];
              muxOutConnector[35] = fifoOut[27][0];
              muxOutConnector[36] = fifoOut[28][0];
              muxOutConnector[37] = fifoOut[29][0];
              muxOutConnector[38] = fifoOut[30][0];
              muxOutConnector[39] = fifoOut[31][0];
              muxOutConnector[40] = fifoOut[32][0];
              muxOutConnector[41] = fifoOut[33][0];
              muxOutConnector[42] = fifoOut[34][0];
              muxOutConnector[43] = fifoOut[35][0];
              muxOutConnector[44] = fifoOut[36][0];
              muxOutConnector[45] = fifoOut[37][0];
              muxOutConnector[46] = fifoOut[38][0];
              muxOutConnector[47] = fifoOut[39][0];
              muxOutConnector[48] = fifoOut[40][0];
              muxOutConnector[49] = fifoOut[41][0];
              muxOutConnector[50] = fifoOut[42][0];
              muxOutConnector[51] = fifoOut[43][0];
       end
       14: begin
              muxOutConnector[0] = fifoOut[49][6];
              muxOutConnector[1] = fifoOut[50][6];
              muxOutConnector[2] = fifoOut[51][6];
              muxOutConnector[3] = fifoOut[26][5];
              muxOutConnector[4] = fifoOut[27][5];
              muxOutConnector[5] = fifoOut[28][5];
              muxOutConnector[6] = fifoOut[29][5];
              muxOutConnector[7] = fifoOut[30][5];
              muxOutConnector[8] = fifoOut[31][5];
              muxOutConnector[9] = fifoOut[32][5];
              muxOutConnector[10] = fifoOut[33][5];
              muxOutConnector[11] = fifoOut[34][5];
              muxOutConnector[12] = fifoOut[35][5];
              muxOutConnector[13] = fifoOut[36][5];
              muxOutConnector[14] = fifoOut[37][5];
              muxOutConnector[15] = fifoOut[38][5];
              muxOutConnector[16] = fifoOut[39][5];
              muxOutConnector[17] = fifoOut[40][5];
              muxOutConnector[18] = fifoOut[41][5];
              muxOutConnector[19] = fifoOut[42][5];
              muxOutConnector[20] = fifoOut[43][5];
              muxOutConnector[21] = fifoOut[44][5];
              muxOutConnector[22] = fifoOut[45][5];
              muxOutConnector[23] = fifoOut[46][5];
              muxOutConnector[24] = fifoOut[47][5];
              muxOutConnector[25] = fifoOut[48][5];
              muxOutConnector[26] = fifoOut[44][1];
              muxOutConnector[27] = fifoOut[45][1];
              muxOutConnector[28] = fifoOut[46][1];
              muxOutConnector[29] = fifoOut[47][1];
              muxOutConnector[30] = fifoOut[48][1];
              muxOutConnector[31] = fifoOut[49][1];
              muxOutConnector[32] = fifoOut[50][1];
              muxOutConnector[33] = fifoOut[51][1];
              muxOutConnector[34] = fifoOut[26][0];
              muxOutConnector[35] = fifoOut[27][0];
              muxOutConnector[36] = fifoOut[28][0];
              muxOutConnector[37] = fifoOut[29][0];
              muxOutConnector[38] = fifoOut[30][0];
              muxOutConnector[39] = fifoOut[31][0];
              muxOutConnector[40] = fifoOut[32][0];
              muxOutConnector[41] = fifoOut[33][0];
              muxOutConnector[42] = fifoOut[34][0];
              muxOutConnector[43] = fifoOut[35][0];
              muxOutConnector[44] = fifoOut[36][0];
              muxOutConnector[45] = fifoOut[37][0];
              muxOutConnector[46] = fifoOut[38][0];
              muxOutConnector[47] = fifoOut[39][0];
              muxOutConnector[48] = fifoOut[40][0];
              muxOutConnector[49] = fifoOut[41][0];
              muxOutConnector[50] = fifoOut[42][0];
              muxOutConnector[51] = fifoOut[43][0];
       end
       15: begin
              muxOutConnector[0] = fifoOut[49][6];
              muxOutConnector[1] = fifoOut[50][6];
              muxOutConnector[2] = fifoOut[51][6];
              muxOutConnector[3] = fifoOut[26][5];
              muxOutConnector[4] = fifoOut[27][5];
              muxOutConnector[5] = fifoOut[28][5];
              muxOutConnector[6] = fifoOut[29][5];
              muxOutConnector[7] = fifoOut[30][5];
              muxOutConnector[8] = fifoOut[31][5];
              muxOutConnector[9] = fifoOut[32][5];
              muxOutConnector[10] = fifoOut[33][5];
              muxOutConnector[11] = fifoOut[34][5];
              muxOutConnector[12] = fifoOut[35][5];
              muxOutConnector[13] = fifoOut[36][5];
              muxOutConnector[14] = fifoOut[37][5];
              muxOutConnector[15] = fifoOut[38][5];
              muxOutConnector[16] = fifoOut[39][5];
              muxOutConnector[17] = fifoOut[40][5];
              muxOutConnector[18] = fifoOut[41][5];
              muxOutConnector[19] = fifoOut[42][5];
              muxOutConnector[20] = fifoOut[43][5];
              muxOutConnector[21] = fifoOut[44][5];
              muxOutConnector[22] = fifoOut[45][5];
              muxOutConnector[23] = fifoOut[46][5];
              muxOutConnector[24] = fifoOut[47][5];
              muxOutConnector[25] = fifoOut[48][5];
              muxOutConnector[26] = fifoOut[44][1];
              muxOutConnector[27] = fifoOut[45][1];
              muxOutConnector[28] = fifoOut[46][1];
              muxOutConnector[29] = fifoOut[47][1];
              muxOutConnector[30] = fifoOut[48][1];
              muxOutConnector[31] = fifoOut[49][1];
              muxOutConnector[32] = fifoOut[50][1];
              muxOutConnector[33] = fifoOut[51][1];
              muxOutConnector[34] = fifoOut[26][0];
              muxOutConnector[35] = fifoOut[27][0];
              muxOutConnector[36] = fifoOut[28][0];
              muxOutConnector[37] = fifoOut[29][0];
              muxOutConnector[38] = fifoOut[30][0];
              muxOutConnector[39] = fifoOut[31][0];
              muxOutConnector[40] = fifoOut[32][0];
              muxOutConnector[41] = fifoOut[33][0];
              muxOutConnector[42] = fifoOut[34][0];
              muxOutConnector[43] = fifoOut[35][0];
              muxOutConnector[44] = fifoOut[36][0];
              muxOutConnector[45] = fifoOut[37][0];
              muxOutConnector[46] = fifoOut[38][0];
              muxOutConnector[47] = fifoOut[39][0];
              muxOutConnector[48] = fifoOut[40][0];
              muxOutConnector[49] = fifoOut[41][0];
              muxOutConnector[50] = fifoOut[42][0];
              muxOutConnector[51] = fifoOut[43][0];
       end
       16: begin
              muxOutConnector[0] = fifoOut[49][6];
              muxOutConnector[1] = fifoOut[50][6];
              muxOutConnector[2] = fifoOut[51][6];
              muxOutConnector[3] = fifoOut[26][5];
              muxOutConnector[4] = fifoOut[27][5];
              muxOutConnector[5] = fifoOut[28][5];
              muxOutConnector[6] = fifoOut[29][5];
              muxOutConnector[7] = fifoOut[30][5];
              muxOutConnector[8] = fifoOut[31][5];
              muxOutConnector[9] = fifoOut[32][5];
              muxOutConnector[10] = fifoOut[33][5];
              muxOutConnector[11] = fifoOut[34][5];
              muxOutConnector[12] = fifoOut[35][5];
              muxOutConnector[13] = fifoOut[36][5];
              muxOutConnector[14] = fifoOut[37][5];
              muxOutConnector[15] = fifoOut[38][5];
              muxOutConnector[16] = fifoOut[39][5];
              muxOutConnector[17] = fifoOut[40][5];
              muxOutConnector[18] = fifoOut[41][5];
              muxOutConnector[19] = fifoOut[42][5];
              muxOutConnector[20] = fifoOut[18][4];
              muxOutConnector[21] = fifoOut[19][4];
              muxOutConnector[22] = fifoOut[20][4];
              muxOutConnector[23] = fifoOut[21][4];
              muxOutConnector[24] = fifoOut[22][4];
              muxOutConnector[25] = fifoOut[23][4];
              muxOutConnector[26] = fifoOut[44][1];
              muxOutConnector[27] = fifoOut[45][1];
              muxOutConnector[28] = fifoOut[46][1];
              muxOutConnector[29] = fifoOut[47][1];
              muxOutConnector[30] = fifoOut[48][1];
              muxOutConnector[31] = fifoOut[49][1];
              muxOutConnector[32] = fifoOut[50][1];
              muxOutConnector[33] = fifoOut[51][1];
              muxOutConnector[34] = fifoOut[26][0];
              muxOutConnector[35] = fifoOut[27][0];
              muxOutConnector[36] = fifoOut[28][0];
              muxOutConnector[37] = fifoOut[29][0];
              muxOutConnector[38] = fifoOut[30][0];
              muxOutConnector[39] = fifoOut[31][0];
              muxOutConnector[40] = fifoOut[32][0];
              muxOutConnector[41] = fifoOut[33][0];
              muxOutConnector[42] = fifoOut[34][0];
              muxOutConnector[43] = fifoOut[35][0];
              muxOutConnector[44] = fifoOut[36][0];
              muxOutConnector[45] = fifoOut[37][0];
              muxOutConnector[46] = fifoOut[38][0];
              muxOutConnector[47] = fifoOut[39][0];
              muxOutConnector[48] = fifoOut[40][0];
              muxOutConnector[49] = fifoOut[41][0];
              muxOutConnector[50] = fifoOut[42][0];
              muxOutConnector[51] = fifoOut[43][0];
       end
       17: begin
              muxOutConnector[0] = fifoOut[24][5];
              muxOutConnector[1] = fifoOut[25][5];
              muxOutConnector[2] = fifoOut[0][4];
              muxOutConnector[3] = fifoOut[1][4];
              muxOutConnector[4] = fifoOut[2][4];
              muxOutConnector[5] = fifoOut[3][4];
              muxOutConnector[6] = fifoOut[4][4];
              muxOutConnector[7] = fifoOut[5][4];
              muxOutConnector[8] = fifoOut[6][4];
              muxOutConnector[9] = fifoOut[7][4];
              muxOutConnector[10] = fifoOut[8][4];
              muxOutConnector[11] = fifoOut[9][4];
              muxOutConnector[12] = fifoOut[10][4];
              muxOutConnector[13] = fifoOut[11][4];
              muxOutConnector[14] = fifoOut[12][4];
              muxOutConnector[15] = fifoOut[13][4];
              muxOutConnector[16] = fifoOut[14][4];
              muxOutConnector[17] = fifoOut[15][4];
              muxOutConnector[18] = fifoOut[16][4];
              muxOutConnector[19] = fifoOut[17][4];
              muxOutConnector[20] = fifoOut[18][4];
              muxOutConnector[21] = fifoOut[19][4];
              muxOutConnector[22] = fifoOut[20][4];
              muxOutConnector[23] = fifoOut[21][4];
              muxOutConnector[24] = fifoOut[22][4];
              muxOutConnector[25] = fifoOut[23][4];
              muxOutConnector[26] = fifoOut[44][1];
              muxOutConnector[27] = fifoOut[45][1];
              muxOutConnector[28] = fifoOut[46][1];
              muxOutConnector[29] = fifoOut[47][1];
              muxOutConnector[30] = fifoOut[48][1];
              muxOutConnector[31] = fifoOut[49][1];
              muxOutConnector[32] = fifoOut[50][1];
              muxOutConnector[33] = fifoOut[51][1];
              muxOutConnector[34] = fifoOut[26][0];
              muxOutConnector[35] = fifoOut[27][0];
              muxOutConnector[36] = fifoOut[28][0];
              muxOutConnector[37] = fifoOut[29][0];
              muxOutConnector[38] = fifoOut[30][0];
              muxOutConnector[39] = fifoOut[31][0];
              muxOutConnector[40] = fifoOut[32][0];
              muxOutConnector[41] = fifoOut[33][0];
              muxOutConnector[42] = fifoOut[34][0];
              muxOutConnector[43] = fifoOut[35][0];
              muxOutConnector[44] = fifoOut[36][0];
              muxOutConnector[45] = fifoOut[37][0];
              muxOutConnector[46] = fifoOut[38][0];
              muxOutConnector[47] = fifoOut[39][0];
              muxOutConnector[48] = fifoOut[40][0];
              muxOutConnector[49] = fifoOut[41][0];
              muxOutConnector[50] = fifoOut[42][0];
              muxOutConnector[51] = fifoOut[43][0];
       end
       18: begin
              muxOutConnector[0] = fifoOut[24][5];
              muxOutConnector[1] = fifoOut[25][5];
              muxOutConnector[2] = fifoOut[0][4];
              muxOutConnector[3] = fifoOut[1][4];
              muxOutConnector[4] = fifoOut[2][4];
              muxOutConnector[5] = fifoOut[3][4];
              muxOutConnector[6] = fifoOut[4][4];
              muxOutConnector[7] = fifoOut[5][4];
              muxOutConnector[8] = fifoOut[6][4];
              muxOutConnector[9] = fifoOut[7][4];
              muxOutConnector[10] = fifoOut[8][4];
              muxOutConnector[11] = fifoOut[9][4];
              muxOutConnector[12] = fifoOut[10][4];
              muxOutConnector[13] = fifoOut[11][4];
              muxOutConnector[14] = fifoOut[12][4];
              muxOutConnector[15] = fifoOut[13][4];
              muxOutConnector[16] = fifoOut[14][4];
              muxOutConnector[17] = fifoOut[15][4];
              muxOutConnector[18] = fifoOut[16][4];
              muxOutConnector[19] = fifoOut[17][4];
              muxOutConnector[20] = fifoOut[18][4];
              muxOutConnector[21] = fifoOut[19][4];
              muxOutConnector[22] = fifoOut[20][4];
              muxOutConnector[23] = fifoOut[21][4];
              muxOutConnector[24] = fifoOut[22][4];
              muxOutConnector[25] = fifoOut[23][4];
              muxOutConnector[26] = fifoOut[44][1];
              muxOutConnector[27] = fifoOut[45][1];
              muxOutConnector[28] = fifoOut[46][1];
              muxOutConnector[29] = fifoOut[47][1];
              muxOutConnector[30] = fifoOut[48][1];
              muxOutConnector[31] = fifoOut[49][1];
              muxOutConnector[32] = fifoOut[50][1];
              muxOutConnector[33] = fifoOut[51][1];
              muxOutConnector[34] = fifoOut[26][0];
              muxOutConnector[35] = fifoOut[27][0];
              muxOutConnector[36] = fifoOut[28][0];
              muxOutConnector[37] = fifoOut[29][0];
              muxOutConnector[38] = fifoOut[30][0];
              muxOutConnector[39] = fifoOut[31][0];
              muxOutConnector[40] = fifoOut[32][0];
              muxOutConnector[41] = fifoOut[33][0];
              muxOutConnector[42] = fifoOut[34][0];
              muxOutConnector[43] = fifoOut[35][0];
              muxOutConnector[44] = fifoOut[36][0];
              muxOutConnector[45] = fifoOut[37][0];
              muxOutConnector[46] = fifoOut[38][0];
              muxOutConnector[47] = fifoOut[39][0];
              muxOutConnector[48] = fifoOut[40][0];
              muxOutConnector[49] = fifoOut[41][0];
              muxOutConnector[50] = fifoOut[42][0];
              muxOutConnector[51] = fifoOut[43][0];
       end
       19: begin
              muxOutConnector[0] = fifoOut[24][5];
              muxOutConnector[1] = fifoOut[25][5];
              muxOutConnector[2] = fifoOut[0][4];
              muxOutConnector[3] = fifoOut[1][4];
              muxOutConnector[4] = fifoOut[2][4];
              muxOutConnector[5] = fifoOut[3][4];
              muxOutConnector[6] = fifoOut[4][4];
              muxOutConnector[7] = fifoOut[5][4];
              muxOutConnector[8] = fifoOut[6][4];
              muxOutConnector[9] = fifoOut[7][4];
              muxOutConnector[10] = fifoOut[8][4];
              muxOutConnector[11] = fifoOut[9][4];
              muxOutConnector[12] = fifoOut[10][4];
              muxOutConnector[13] = fifoOut[11][4];
              muxOutConnector[14] = fifoOut[12][4];
              muxOutConnector[15] = fifoOut[13][4];
              muxOutConnector[16] = fifoOut[14][4];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[44][1];
              muxOutConnector[27] = fifoOut[45][1];
              muxOutConnector[28] = fifoOut[46][1];
              muxOutConnector[29] = fifoOut[47][1];
              muxOutConnector[30] = fifoOut[48][1];
              muxOutConnector[31] = fifoOut[49][1];
              muxOutConnector[32] = fifoOut[50][1];
              muxOutConnector[33] = fifoOut[51][1];
              muxOutConnector[34] = fifoOut[26][0];
              muxOutConnector[35] = fifoOut[27][0];
              muxOutConnector[36] = fifoOut[28][0];
              muxOutConnector[37] = fifoOut[29][0];
              muxOutConnector[38] = fifoOut[30][0];
              muxOutConnector[39] = fifoOut[31][0];
              muxOutConnector[40] = fifoOut[32][0];
              muxOutConnector[41] = fifoOut[33][0];
              muxOutConnector[42] = fifoOut[34][0];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
