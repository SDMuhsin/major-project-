`timescale 1ns / 1ps
module LMem0To1_511_circ7_ys_scripted(
        muxOut,
        ly0In,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 14;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

reg   feedback_en;
reg [ w - 1 : 0 ]column_1[ r - 1 : 0 ];
reg chip_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(chip_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= column_1[i];
         end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
  feedback_en=rd_en;
      if(wr_en)begin
        chip_en=wr_en;
      end
      else begin
        chip_en=feedback_en;
      end
   if(feedback_en)begin
      for(i = r-1; i > -1; i=i-1) begin
        column_1[i] <= fifoOut[i][c-1];
      end
   end
   else begin
      for(i = r-1; i > -1; i=i-1) begin
        column_1[i] <= ly0InConnector[i];
      end
    end
end
always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[2][12];
              muxOutConnector[1] = fifoOut[3][12];
              muxOutConnector[2] = fifoOut[4][12];
              muxOutConnector[3] = fifoOut[5][12];
              muxOutConnector[4] = fifoOut[6][12];
              muxOutConnector[5] = fifoOut[7][12];
              muxOutConnector[6] = fifoOut[8][12];
              muxOutConnector[7] = fifoOut[9][12];
              muxOutConnector[8] = fifoOut[10][12];
              muxOutConnector[9] = fifoOut[11][12];
              muxOutConnector[10] = fifoOut[12][12];
              muxOutConnector[11] = fifoOut[13][12];
              muxOutConnector[12] = fifoOut[14][12];
              muxOutConnector[13] = fifoOut[15][12];
              muxOutConnector[14] = fifoOut[16][12];
              muxOutConnector[15] = fifoOut[17][12];
              muxOutConnector[16] = fifoOut[18][12];
              muxOutConnector[17] = fifoOut[19][12];
              muxOutConnector[18] = fifoOut[20][12];
              muxOutConnector[19] = fifoOut[21][12];
              muxOutConnector[20] = fifoOut[22][12];
              muxOutConnector[21] = fifoOut[23][12];
              muxOutConnector[22] = fifoOut[24][12];
              muxOutConnector[23] = fifoOut[25][12];
              muxOutConnector[24] = fifoOut[0][11];
              muxOutConnector[25] = fifoOut[1][11];
              muxOutConnector[26] = fifoOut[20][3];
              muxOutConnector[27] = fifoOut[21][3];
              muxOutConnector[28] = fifoOut[22][3];
              muxOutConnector[29] = fifoOut[23][3];
              muxOutConnector[30] = fifoOut[24][3];
              muxOutConnector[31] = fifoOut[25][3];
              muxOutConnector[32] = fifoOut[0][2];
              muxOutConnector[33] = fifoOut[1][2];
              muxOutConnector[34] = fifoOut[2][2];
              muxOutConnector[35] = fifoOut[3][2];
              muxOutConnector[36] = fifoOut[4][2];
              muxOutConnector[37] = fifoOut[5][2];
              muxOutConnector[38] = fifoOut[6][2];
              muxOutConnector[39] = fifoOut[7][2];
              muxOutConnector[40] = fifoOut[8][2];
              muxOutConnector[41] = fifoOut[9][2];
              muxOutConnector[42] = fifoOut[10][2];
              muxOutConnector[43] = fifoOut[11][2];
              muxOutConnector[44] = fifoOut[12][2];
              muxOutConnector[45] = fifoOut[13][2];
              muxOutConnector[46] = fifoOut[14][2];
              muxOutConnector[47] = fifoOut[15][2];
              muxOutConnector[48] = fifoOut[16][2];
              muxOutConnector[49] = fifoOut[17][2];
              muxOutConnector[50] = fifoOut[18][2];
              muxOutConnector[51] = fifoOut[19][2];
       end
       1: begin
              muxOutConnector[0] = fifoOut[2][12];
              muxOutConnector[1] = fifoOut[3][12];
              muxOutConnector[2] = fifoOut[4][12];
              muxOutConnector[3] = fifoOut[5][12];
              muxOutConnector[4] = fifoOut[6][12];
              muxOutConnector[5] = fifoOut[7][12];
              muxOutConnector[6] = fifoOut[8][12];
              muxOutConnector[7] = fifoOut[9][12];
              muxOutConnector[8] = fifoOut[10][12];
              muxOutConnector[9] = fifoOut[11][12];
              muxOutConnector[10] = fifoOut[12][12];
              muxOutConnector[11] = fifoOut[13][12];
              muxOutConnector[12] = fifoOut[14][12];
              muxOutConnector[13] = fifoOut[15][12];
              muxOutConnector[14] = fifoOut[16][12];
              muxOutConnector[15] = fifoOut[17][12];
              muxOutConnector[16] = fifoOut[18][12];
              muxOutConnector[17] = fifoOut[19][12];
              muxOutConnector[18] = fifoOut[20][12];
              muxOutConnector[19] = fifoOut[21][12];
              muxOutConnector[20] = fifoOut[22][12];
              muxOutConnector[21] = fifoOut[23][12];
              muxOutConnector[22] = fifoOut[24][12];
              muxOutConnector[23] = fifoOut[25][12];
              muxOutConnector[24] = fifoOut[0][11];
              muxOutConnector[25] = fifoOut[1][11];
              muxOutConnector[26] = fifoOut[20][3];
              muxOutConnector[27] = fifoOut[21][3];
              muxOutConnector[28] = fifoOut[22][3];
              muxOutConnector[29] = fifoOut[23][3];
              muxOutConnector[30] = fifoOut[24][3];
              muxOutConnector[31] = fifoOut[25][3];
              muxOutConnector[32] = fifoOut[0][2];
              muxOutConnector[33] = fifoOut[1][2];
              muxOutConnector[34] = fifoOut[2][2];
              muxOutConnector[35] = fifoOut[3][2];
              muxOutConnector[36] = fifoOut[4][2];
              muxOutConnector[37] = fifoOut[5][2];
              muxOutConnector[38] = fifoOut[6][2];
              muxOutConnector[39] = fifoOut[7][2];
              muxOutConnector[40] = fifoOut[8][2];
              muxOutConnector[41] = fifoOut[9][2];
              muxOutConnector[42] = fifoOut[10][2];
              muxOutConnector[43] = fifoOut[11][2];
              muxOutConnector[44] = fifoOut[12][2];
              muxOutConnector[45] = fifoOut[13][2];
              muxOutConnector[46] = fifoOut[14][2];
              muxOutConnector[47] = fifoOut[15][2];
              muxOutConnector[48] = fifoOut[16][2];
              muxOutConnector[49] = fifoOut[17][2];
              muxOutConnector[50] = fifoOut[18][2];
              muxOutConnector[51] = fifoOut[19][2];
       end
       2: begin
              muxOutConnector[0] = fifoOut[2][12];
              muxOutConnector[1] = fifoOut[3][12];
              muxOutConnector[2] = fifoOut[4][12];
              muxOutConnector[3] = fifoOut[5][12];
              muxOutConnector[4] = fifoOut[6][12];
              muxOutConnector[5] = fifoOut[7][12];
              muxOutConnector[6] = fifoOut[8][12];
              muxOutConnector[7] = fifoOut[9][12];
              muxOutConnector[8] = fifoOut[10][12];
              muxOutConnector[9] = fifoOut[11][12];
              muxOutConnector[10] = fifoOut[12][12];
              muxOutConnector[11] = fifoOut[13][12];
              muxOutConnector[12] = fifoOut[14][12];
              muxOutConnector[13] = fifoOut[15][12];
              muxOutConnector[14] = fifoOut[16][12];
              muxOutConnector[15] = fifoOut[17][12];
              muxOutConnector[16] = fifoOut[18][12];
              muxOutConnector[17] = fifoOut[19][12];
              muxOutConnector[18] = fifoOut[20][12];
              muxOutConnector[19] = fifoOut[21][12];
              muxOutConnector[20] = fifoOut[22][12];
              muxOutConnector[21] = fifoOut[23][12];
              muxOutConnector[22] = fifoOut[24][12];
              muxOutConnector[23] = fifoOut[25][12];
              muxOutConnector[24] = fifoOut[0][11];
              muxOutConnector[25] = fifoOut[1][11];
              muxOutConnector[26] = fifoOut[20][3];
              muxOutConnector[27] = fifoOut[21][3];
              muxOutConnector[28] = fifoOut[22][3];
              muxOutConnector[29] = fifoOut[23][3];
              muxOutConnector[30] = fifoOut[24][3];
              muxOutConnector[31] = fifoOut[25][3];
              muxOutConnector[32] = fifoOut[0][2];
              muxOutConnector[33] = fifoOut[1][2];
              muxOutConnector[34] = fifoOut[2][2];
              muxOutConnector[35] = fifoOut[3][2];
              muxOutConnector[36] = fifoOut[4][2];
              muxOutConnector[37] = fifoOut[5][2];
              muxOutConnector[38] = fifoOut[6][2];
              muxOutConnector[39] = fifoOut[7][2];
              muxOutConnector[40] = fifoOut[8][2];
              muxOutConnector[41] = fifoOut[9][2];
              muxOutConnector[42] = fifoOut[10][2];
              muxOutConnector[43] = fifoOut[11][2];
              muxOutConnector[44] = fifoOut[12][2];
              muxOutConnector[45] = fifoOut[13][2];
              muxOutConnector[46] = fifoOut[14][2];
              muxOutConnector[47] = fifoOut[15][2];
              muxOutConnector[48] = fifoOut[16][2];
              muxOutConnector[49] = fifoOut[31][1];
              muxOutConnector[50] = fifoOut[32][1];
              muxOutConnector[51] = fifoOut[33][1];
       end
       3: begin
              muxOutConnector[0] = fifoOut[2][12];
              muxOutConnector[1] = fifoOut[3][12];
              muxOutConnector[2] = fifoOut[4][12];
              muxOutConnector[3] = fifoOut[5][12];
              muxOutConnector[4] = fifoOut[6][12];
              muxOutConnector[5] = fifoOut[7][12];
              muxOutConnector[6] = fifoOut[8][12];
              muxOutConnector[7] = fifoOut[9][12];
              muxOutConnector[8] = fifoOut[10][12];
              muxOutConnector[9] = fifoOut[11][12];
              muxOutConnector[10] = fifoOut[12][12];
              muxOutConnector[11] = fifoOut[13][12];
              muxOutConnector[12] = fifoOut[14][12];
              muxOutConnector[13] = fifoOut[15][12];
              muxOutConnector[14] = fifoOut[16][12];
              muxOutConnector[15] = fifoOut[17][12];
              muxOutConnector[16] = fifoOut[18][12];
              muxOutConnector[17] = fifoOut[19][12];
              muxOutConnector[18] = fifoOut[20][12];
              muxOutConnector[19] = fifoOut[21][12];
              muxOutConnector[20] = fifoOut[22][12];
              muxOutConnector[21] = fifoOut[23][12];
              muxOutConnector[22] = fifoOut[24][12];
              muxOutConnector[23] = fifoOut[25][12];
              muxOutConnector[24] = fifoOut[0][11];
              muxOutConnector[25] = fifoOut[1][11];
              muxOutConnector[26] = fifoOut[34][2];
              muxOutConnector[27] = fifoOut[35][2];
              muxOutConnector[28] = fifoOut[36][2];
              muxOutConnector[29] = fifoOut[37][2];
              muxOutConnector[30] = fifoOut[38][2];
              muxOutConnector[31] = fifoOut[39][2];
              muxOutConnector[32] = fifoOut[40][2];
              muxOutConnector[33] = fifoOut[41][2];
              muxOutConnector[34] = fifoOut[42][2];
              muxOutConnector[35] = fifoOut[43][2];
              muxOutConnector[36] = fifoOut[44][2];
              muxOutConnector[37] = fifoOut[45][2];
              muxOutConnector[38] = fifoOut[46][2];
              muxOutConnector[39] = fifoOut[47][2];
              muxOutConnector[40] = fifoOut[48][2];
              muxOutConnector[41] = fifoOut[49][2];
              muxOutConnector[42] = fifoOut[50][2];
              muxOutConnector[43] = fifoOut[51][2];
              muxOutConnector[44] = fifoOut[26][1];
              muxOutConnector[45] = fifoOut[27][1];
              muxOutConnector[46] = fifoOut[28][1];
              muxOutConnector[47] = fifoOut[29][1];
              muxOutConnector[48] = fifoOut[30][1];
              muxOutConnector[49] = fifoOut[31][1];
              muxOutConnector[50] = fifoOut[32][1];
              muxOutConnector[51] = fifoOut[33][1];
       end
       4: begin
              muxOutConnector[0] = fifoOut[2][12];
              muxOutConnector[1] = fifoOut[3][12];
              muxOutConnector[2] = fifoOut[4][12];
              muxOutConnector[3] = fifoOut[5][12];
              muxOutConnector[4] = fifoOut[6][12];
              muxOutConnector[5] = fifoOut[7][12];
              muxOutConnector[6] = fifoOut[8][12];
              muxOutConnector[7] = fifoOut[9][12];
              muxOutConnector[8] = fifoOut[10][12];
              muxOutConnector[9] = fifoOut[11][12];
              muxOutConnector[10] = fifoOut[12][12];
              muxOutConnector[11] = fifoOut[13][12];
              muxOutConnector[12] = fifoOut[14][12];
              muxOutConnector[13] = fifoOut[15][12];
              muxOutConnector[14] = fifoOut[16][12];
              muxOutConnector[15] = fifoOut[17][12];
              muxOutConnector[16] = fifoOut[18][12];
              muxOutConnector[17] = fifoOut[19][12];
              muxOutConnector[18] = fifoOut[20][12];
              muxOutConnector[19] = fifoOut[21][12];
              muxOutConnector[20] = fifoOut[22][12];
              muxOutConnector[21] = fifoOut[23][12];
              muxOutConnector[22] = fifoOut[24][12];
              muxOutConnector[23] = fifoOut[25][12];
              muxOutConnector[24] = fifoOut[0][11];
              muxOutConnector[25] = fifoOut[1][11];
              muxOutConnector[26] = fifoOut[34][2];
              muxOutConnector[27] = fifoOut[35][2];
              muxOutConnector[28] = fifoOut[36][2];
              muxOutConnector[29] = fifoOut[37][2];
              muxOutConnector[30] = fifoOut[38][2];
              muxOutConnector[31] = fifoOut[39][2];
              muxOutConnector[32] = fifoOut[40][2];
              muxOutConnector[33] = fifoOut[41][2];
              muxOutConnector[34] = fifoOut[42][2];
              muxOutConnector[35] = fifoOut[43][2];
              muxOutConnector[36] = fifoOut[44][2];
              muxOutConnector[37] = fifoOut[45][2];
              muxOutConnector[38] = fifoOut[46][2];
              muxOutConnector[39] = fifoOut[47][2];
              muxOutConnector[40] = fifoOut[48][2];
              muxOutConnector[41] = fifoOut[49][2];
              muxOutConnector[42] = fifoOut[50][2];
              muxOutConnector[43] = fifoOut[51][2];
              muxOutConnector[44] = fifoOut[26][1];
              muxOutConnector[45] = fifoOut[27][1];
              muxOutConnector[46] = fifoOut[28][1];
              muxOutConnector[47] = fifoOut[29][1];
              muxOutConnector[48] = fifoOut[30][1];
              muxOutConnector[49] = fifoOut[31][1];
              muxOutConnector[50] = fifoOut[32][1];
              muxOutConnector[51] = fifoOut[33][1];
       end
       5: begin
              muxOutConnector[0] = fifoOut[2][12];
              muxOutConnector[1] = fifoOut[3][12];
              muxOutConnector[2] = fifoOut[4][12];
              muxOutConnector[3] = fifoOut[5][12];
              muxOutConnector[4] = fifoOut[6][12];
              muxOutConnector[5] = fifoOut[7][12];
              muxOutConnector[6] = fifoOut[8][12];
              muxOutConnector[7] = fifoOut[9][12];
              muxOutConnector[8] = fifoOut[10][12];
              muxOutConnector[9] = fifoOut[11][12];
              muxOutConnector[10] = fifoOut[12][12];
              muxOutConnector[11] = fifoOut[13][12];
              muxOutConnector[12] = fifoOut[14][12];
              muxOutConnector[13] = fifoOut[15][12];
              muxOutConnector[14] = fifoOut[16][12];
              muxOutConnector[15] = fifoOut[17][12];
              muxOutConnector[16] = fifoOut[18][12];
              muxOutConnector[17] = fifoOut[19][12];
              muxOutConnector[18] = fifoOut[20][12];
              muxOutConnector[19] = fifoOut[21][12];
              muxOutConnector[20] = fifoOut[22][12];
              muxOutConnector[21] = fifoOut[23][12];
              muxOutConnector[22] = fifoOut[24][12];
              muxOutConnector[23] = fifoOut[25][12];
              muxOutConnector[24] = fifoOut[0][11];
              muxOutConnector[25] = fifoOut[1][11];
              muxOutConnector[26] = fifoOut[34][2];
              muxOutConnector[27] = fifoOut[35][2];
              muxOutConnector[28] = fifoOut[36][2];
              muxOutConnector[29] = fifoOut[37][2];
              muxOutConnector[30] = fifoOut[38][2];
              muxOutConnector[31] = fifoOut[39][2];
              muxOutConnector[32] = fifoOut[40][2];
              muxOutConnector[33] = fifoOut[41][2];
              muxOutConnector[34] = fifoOut[42][2];
              muxOutConnector[35] = fifoOut[43][2];
              muxOutConnector[36] = fifoOut[44][2];
              muxOutConnector[37] = fifoOut[45][2];
              muxOutConnector[38] = fifoOut[46][2];
              muxOutConnector[39] = fifoOut[47][2];
              muxOutConnector[40] = fifoOut[48][2];
              muxOutConnector[41] = fifoOut[49][2];
              muxOutConnector[42] = fifoOut[50][2];
              muxOutConnector[43] = fifoOut[51][2];
              muxOutConnector[44] = fifoOut[26][1];
              muxOutConnector[45] = fifoOut[27][1];
              muxOutConnector[46] = fifoOut[28][1];
              muxOutConnector[47] = fifoOut[29][1];
              muxOutConnector[48] = fifoOut[30][1];
              muxOutConnector[49] = fifoOut[31][1];
              muxOutConnector[50] = fifoOut[32][1];
              muxOutConnector[51] = fifoOut[33][1];
       end
       6: begin
              muxOutConnector[0] = fifoOut[2][12];
              muxOutConnector[1] = fifoOut[3][12];
              muxOutConnector[2] = fifoOut[4][12];
              muxOutConnector[3] = fifoOut[5][12];
              muxOutConnector[4] = fifoOut[6][12];
              muxOutConnector[5] = fifoOut[7][12];
              muxOutConnector[6] = fifoOut[8][12];
              muxOutConnector[7] = fifoOut[9][12];
              muxOutConnector[8] = fifoOut[10][12];
              muxOutConnector[9] = fifoOut[11][12];
              muxOutConnector[10] = fifoOut[12][12];
              muxOutConnector[11] = fifoOut[13][12];
              muxOutConnector[12] = fifoOut[14][12];
              muxOutConnector[13] = fifoOut[15][12];
              muxOutConnector[14] = fifoOut[16][12];
              muxOutConnector[15] = fifoOut[17][12];
              muxOutConnector[16] = fifoOut[18][12];
              muxOutConnector[17] = fifoOut[19][12];
              muxOutConnector[18] = fifoOut[20][12];
              muxOutConnector[19] = fifoOut[21][12];
              muxOutConnector[20] = fifoOut[22][12];
              muxOutConnector[21] = fifoOut[23][12];
              muxOutConnector[22] = fifoOut[24][12];
              muxOutConnector[23] = fifoOut[25][12];
              muxOutConnector[24] = fifoOut[0][11];
              muxOutConnector[25] = fifoOut[1][11];
              muxOutConnector[26] = fifoOut[34][2];
              muxOutConnector[27] = fifoOut[35][2];
              muxOutConnector[28] = fifoOut[36][2];
              muxOutConnector[29] = fifoOut[37][2];
              muxOutConnector[30] = fifoOut[38][2];
              muxOutConnector[31] = fifoOut[39][2];
              muxOutConnector[32] = fifoOut[40][2];
              muxOutConnector[33] = fifoOut[41][2];
              muxOutConnector[34] = fifoOut[42][2];
              muxOutConnector[35] = fifoOut[43][2];
              muxOutConnector[36] = fifoOut[44][2];
              muxOutConnector[37] = fifoOut[45][2];
              muxOutConnector[38] = fifoOut[46][2];
              muxOutConnector[39] = fifoOut[47][2];
              muxOutConnector[40] = fifoOut[48][2];
              muxOutConnector[41] = fifoOut[49][2];
              muxOutConnector[42] = fifoOut[50][2];
              muxOutConnector[43] = fifoOut[51][2];
              muxOutConnector[44] = fifoOut[26][1];
              muxOutConnector[45] = fifoOut[27][1];
              muxOutConnector[46] = fifoOut[28][1];
              muxOutConnector[47] = fifoOut[29][1];
              muxOutConnector[48] = fifoOut[30][1];
              muxOutConnector[49] = fifoOut[31][1];
              muxOutConnector[50] = fifoOut[32][1];
              muxOutConnector[51] = fifoOut[33][1];
       end
       7: begin
              muxOutConnector[0] = fifoOut[2][12];
              muxOutConnector[1] = fifoOut[3][12];
              muxOutConnector[2] = fifoOut[4][12];
              muxOutConnector[3] = fifoOut[5][12];
              muxOutConnector[4] = fifoOut[6][12];
              muxOutConnector[5] = fifoOut[7][12];
              muxOutConnector[6] = fifoOut[8][12];
              muxOutConnector[7] = fifoOut[9][12];
              muxOutConnector[8] = fifoOut[10][12];
              muxOutConnector[9] = fifoOut[11][12];
              muxOutConnector[10] = fifoOut[12][12];
              muxOutConnector[11] = fifoOut[13][12];
              muxOutConnector[12] = fifoOut[14][12];
              muxOutConnector[13] = fifoOut[15][12];
              muxOutConnector[14] = fifoOut[16][12];
              muxOutConnector[15] = fifoOut[17][12];
              muxOutConnector[16] = fifoOut[18][12];
              muxOutConnector[17] = fifoOut[19][12];
              muxOutConnector[18] = fifoOut[20][12];
              muxOutConnector[19] = fifoOut[21][12];
              muxOutConnector[20] = fifoOut[22][12];
              muxOutConnector[21] = fifoOut[23][12];
              muxOutConnector[22] = fifoOut[24][12];
              muxOutConnector[23] = fifoOut[25][12];
              muxOutConnector[24] = fifoOut[0][11];
              muxOutConnector[25] = fifoOut[1][11];
              muxOutConnector[26] = fifoOut[34][2];
              muxOutConnector[27] = fifoOut[35][2];
              muxOutConnector[28] = fifoOut[36][2];
              muxOutConnector[29] = fifoOut[37][2];
              muxOutConnector[30] = fifoOut[38][2];
              muxOutConnector[31] = fifoOut[39][2];
              muxOutConnector[32] = fifoOut[40][2];
              muxOutConnector[33] = fifoOut[41][2];
              muxOutConnector[34] = fifoOut[42][2];
              muxOutConnector[35] = fifoOut[43][2];
              muxOutConnector[36] = fifoOut[44][2];
              muxOutConnector[37] = fifoOut[45][2];
              muxOutConnector[38] = fifoOut[46][2];
              muxOutConnector[39] = fifoOut[47][2];
              muxOutConnector[40] = fifoOut[48][2];
              muxOutConnector[41] = fifoOut[49][2];
              muxOutConnector[42] = fifoOut[50][2];
              muxOutConnector[43] = fifoOut[51][2];
              muxOutConnector[44] = fifoOut[26][1];
              muxOutConnector[45] = fifoOut[27][1];
              muxOutConnector[46] = fifoOut[28][1];
              muxOutConnector[47] = fifoOut[29][1];
              muxOutConnector[48] = fifoOut[30][1];
              muxOutConnector[49] = fifoOut[31][1];
              muxOutConnector[50] = fifoOut[32][1];
              muxOutConnector[51] = fifoOut[33][1];
       end
       8: begin
              muxOutConnector[0] = fifoOut[2][12];
              muxOutConnector[1] = fifoOut[3][12];
              muxOutConnector[2] = fifoOut[4][12];
              muxOutConnector[3] = fifoOut[5][12];
              muxOutConnector[4] = fifoOut[6][12];
              muxOutConnector[5] = fifoOut[7][12];
              muxOutConnector[6] = fifoOut[8][12];
              muxOutConnector[7] = fifoOut[9][12];
              muxOutConnector[8] = fifoOut[10][12];
              muxOutConnector[9] = fifoOut[11][12];
              muxOutConnector[10] = fifoOut[12][12];
              muxOutConnector[11] = fifoOut[13][12];
              muxOutConnector[12] = fifoOut[14][12];
              muxOutConnector[13] = fifoOut[15][12];
              muxOutConnector[14] = fifoOut[16][12];
              muxOutConnector[15] = fifoOut[17][12];
              muxOutConnector[16] = fifoOut[18][12];
              muxOutConnector[17] = fifoOut[19][12];
              muxOutConnector[18] = fifoOut[20][12];
              muxOutConnector[19] = fifoOut[21][12];
              muxOutConnector[20] = fifoOut[22][12];
              muxOutConnector[21] = fifoOut[23][12];
              muxOutConnector[22] = fifoOut[24][12];
              muxOutConnector[23] = fifoOut[25][12];
              muxOutConnector[24] = fifoOut[0][11];
              muxOutConnector[25] = fifoOut[1][11];
              muxOutConnector[26] = fifoOut[34][2];
              muxOutConnector[27] = fifoOut[35][2];
              muxOutConnector[28] = fifoOut[36][2];
              muxOutConnector[29] = fifoOut[37][2];
              muxOutConnector[30] = fifoOut[38][2];
              muxOutConnector[31] = fifoOut[39][2];
              muxOutConnector[32] = fifoOut[40][2];
              muxOutConnector[33] = fifoOut[41][2];
              muxOutConnector[34] = fifoOut[42][2];
              muxOutConnector[35] = fifoOut[43][2];
              muxOutConnector[36] = fifoOut[44][2];
              muxOutConnector[37] = fifoOut[45][2];
              muxOutConnector[38] = fifoOut[46][2];
              muxOutConnector[39] = fifoOut[47][2];
              muxOutConnector[40] = fifoOut[48][2];
              muxOutConnector[41] = fifoOut[49][2];
              muxOutConnector[42] = fifoOut[50][2];
              muxOutConnector[43] = fifoOut[51][2];
              muxOutConnector[44] = fifoOut[26][1];
              muxOutConnector[45] = fifoOut[27][1];
              muxOutConnector[46] = fifoOut[28][1];
              muxOutConnector[47] = fifoOut[29][1];
              muxOutConnector[48] = fifoOut[30][1];
              muxOutConnector[49] = fifoOut[0][7];
              muxOutConnector[50] = fifoOut[1][7];
              muxOutConnector[51] = fifoOut[2][7];
       end
       9: begin
              muxOutConnector[0] = fifoOut[2][12];
              muxOutConnector[1] = fifoOut[3][12];
              muxOutConnector[2] = fifoOut[4][12];
              muxOutConnector[3] = fifoOut[5][12];
              muxOutConnector[4] = fifoOut[6][12];
              muxOutConnector[5] = fifoOut[7][12];
              muxOutConnector[6] = fifoOut[8][12];
              muxOutConnector[7] = fifoOut[9][12];
              muxOutConnector[8] = fifoOut[10][12];
              muxOutConnector[9] = fifoOut[11][12];
              muxOutConnector[10] = fifoOut[12][12];
              muxOutConnector[11] = fifoOut[13][12];
              muxOutConnector[12] = fifoOut[14][12];
              muxOutConnector[13] = fifoOut[15][12];
              muxOutConnector[14] = fifoOut[16][12];
              muxOutConnector[15] = fifoOut[17][12];
              muxOutConnector[16] = fifoOut[18][12];
              muxOutConnector[17] = fifoOut[19][12];
              muxOutConnector[18] = fifoOut[20][12];
              muxOutConnector[19] = fifoOut[21][12];
              muxOutConnector[20] = fifoOut[22][12];
              muxOutConnector[21] = fifoOut[23][12];
              muxOutConnector[22] = fifoOut[24][12];
              muxOutConnector[23] = fifoOut[25][12];
              muxOutConnector[24] = fifoOut[0][11];
              muxOutConnector[25] = fifoOut[1][11];
              muxOutConnector[26] = fifoOut[3][8];
              muxOutConnector[27] = fifoOut[4][8];
              muxOutConnector[28] = fifoOut[5][8];
              muxOutConnector[29] = fifoOut[6][8];
              muxOutConnector[30] = fifoOut[7][8];
              muxOutConnector[31] = fifoOut[8][8];
              muxOutConnector[32] = fifoOut[9][8];
              muxOutConnector[33] = fifoOut[10][8];
              muxOutConnector[34] = fifoOut[11][8];
              muxOutConnector[35] = fifoOut[12][8];
              muxOutConnector[36] = fifoOut[13][8];
              muxOutConnector[37] = fifoOut[14][8];
              muxOutConnector[38] = fifoOut[15][8];
              muxOutConnector[39] = fifoOut[16][8];
              muxOutConnector[40] = fifoOut[17][8];
              muxOutConnector[41] = fifoOut[18][8];
              muxOutConnector[42] = fifoOut[19][8];
              muxOutConnector[43] = fifoOut[20][8];
              muxOutConnector[44] = fifoOut[21][8];
              muxOutConnector[45] = fifoOut[22][8];
              muxOutConnector[46] = fifoOut[23][8];
              muxOutConnector[47] = fifoOut[24][8];
              muxOutConnector[48] = fifoOut[25][8];
              muxOutConnector[49] = fifoOut[0][7];
              muxOutConnector[50] = fifoOut[1][7];
              muxOutConnector[51] = fifoOut[2][7];
       end
       10: begin
              muxOutConnector[0] = fifoOut[2][12];
              muxOutConnector[1] = fifoOut[3][12];
              muxOutConnector[2] = fifoOut[4][12];
              muxOutConnector[3] = fifoOut[5][12];
              muxOutConnector[4] = fifoOut[6][12];
              muxOutConnector[5] = fifoOut[7][12];
              muxOutConnector[6] = fifoOut[8][12];
              muxOutConnector[7] = fifoOut[9][12];
              muxOutConnector[8] = fifoOut[10][12];
              muxOutConnector[9] = fifoOut[11][12];
              muxOutConnector[10] = fifoOut[12][12];
              muxOutConnector[11] = fifoOut[13][12];
              muxOutConnector[12] = fifoOut[14][12];
              muxOutConnector[13] = fifoOut[15][12];
              muxOutConnector[14] = fifoOut[16][12];
              muxOutConnector[15] = fifoOut[17][12];
              muxOutConnector[16] = fifoOut[18][12];
              muxOutConnector[17] = fifoOut[19][12];
              muxOutConnector[18] = fifoOut[20][12];
              muxOutConnector[19] = fifoOut[21][12];
              muxOutConnector[20] = fifoOut[22][12];
              muxOutConnector[21] = fifoOut[23][12];
              muxOutConnector[22] = fifoOut[24][12];
              muxOutConnector[23] = fifoOut[25][12];
              muxOutConnector[24] = fifoOut[0][11];
              muxOutConnector[25] = fifoOut[1][11];
              muxOutConnector[26] = fifoOut[3][8];
              muxOutConnector[27] = fifoOut[4][8];
              muxOutConnector[28] = fifoOut[5][8];
              muxOutConnector[29] = fifoOut[6][8];
              muxOutConnector[30] = fifoOut[7][8];
              muxOutConnector[31] = fifoOut[8][8];
              muxOutConnector[32] = fifoOut[9][8];
              muxOutConnector[33] = fifoOut[10][8];
              muxOutConnector[34] = fifoOut[11][8];
              muxOutConnector[35] = fifoOut[12][8];
              muxOutConnector[36] = fifoOut[13][8];
              muxOutConnector[37] = fifoOut[14][8];
              muxOutConnector[38] = fifoOut[15][8];
              muxOutConnector[39] = fifoOut[16][8];
              muxOutConnector[40] = fifoOut[17][8];
              muxOutConnector[41] = fifoOut[18][8];
              muxOutConnector[42] = fifoOut[19][8];
              muxOutConnector[43] = fifoOut[20][8];
              muxOutConnector[44] = fifoOut[21][8];
              muxOutConnector[45] = fifoOut[22][8];
              muxOutConnector[46] = fifoOut[23][8];
              muxOutConnector[47] = fifoOut[24][8];
              muxOutConnector[48] = fifoOut[25][8];
              muxOutConnector[49] = fifoOut[0][7];
              muxOutConnector[50] = fifoOut[1][7];
              muxOutConnector[51] = fifoOut[2][7];
       end
       11: begin
              muxOutConnector[0] = fifoOut[2][12];
              muxOutConnector[1] = fifoOut[3][12];
              muxOutConnector[2] = fifoOut[4][12];
              muxOutConnector[3] = fifoOut[5][12];
              muxOutConnector[4] = fifoOut[6][12];
              muxOutConnector[5] = fifoOut[7][12];
              muxOutConnector[6] = fifoOut[8][12];
              muxOutConnector[7] = fifoOut[9][12];
              muxOutConnector[8] = fifoOut[10][12];
              muxOutConnector[9] = fifoOut[11][12];
              muxOutConnector[10] = fifoOut[12][12];
              muxOutConnector[11] = fifoOut[13][12];
              muxOutConnector[12] = fifoOut[14][12];
              muxOutConnector[13] = fifoOut[15][12];
              muxOutConnector[14] = fifoOut[16][12];
              muxOutConnector[15] = fifoOut[17][12];
              muxOutConnector[16] = fifoOut[18][12];
              muxOutConnector[17] = fifoOut[19][12];
              muxOutConnector[18] = fifoOut[20][12];
              muxOutConnector[19] = fifoOut[21][12];
              muxOutConnector[20] = fifoOut[22][12];
              muxOutConnector[21] = fifoOut[23][12];
              muxOutConnector[22] = fifoOut[24][12];
              muxOutConnector[23] = fifoOut[25][12];
              muxOutConnector[24] = fifoOut[0][11];
              muxOutConnector[25] = fifoOut[1][11];
              muxOutConnector[26] = fifoOut[3][8];
              muxOutConnector[27] = fifoOut[4][8];
              muxOutConnector[28] = fifoOut[5][8];
              muxOutConnector[29] = fifoOut[6][8];
              muxOutConnector[30] = fifoOut[7][8];
              muxOutConnector[31] = fifoOut[8][8];
              muxOutConnector[32] = fifoOut[9][8];
              muxOutConnector[33] = fifoOut[10][8];
              muxOutConnector[34] = fifoOut[11][8];
              muxOutConnector[35] = fifoOut[12][8];
              muxOutConnector[36] = fifoOut[13][8];
              muxOutConnector[37] = fifoOut[14][8];
              muxOutConnector[38] = fifoOut[15][8];
              muxOutConnector[39] = fifoOut[16][8];
              muxOutConnector[40] = fifoOut[17][8];
              muxOutConnector[41] = fifoOut[18][8];
              muxOutConnector[42] = fifoOut[19][8];
              muxOutConnector[43] = fifoOut[20][8];
              muxOutConnector[44] = fifoOut[21][8];
              muxOutConnector[45] = fifoOut[22][8];
              muxOutConnector[46] = fifoOut[23][8];
              muxOutConnector[47] = fifoOut[24][8];
              muxOutConnector[48] = fifoOut[25][8];
              muxOutConnector[49] = fifoOut[0][7];
              muxOutConnector[50] = fifoOut[1][7];
              muxOutConnector[51] = fifoOut[2][7];
       end
       12: begin
              muxOutConnector[0] = fifoOut[2][12];
              muxOutConnector[1] = fifoOut[3][12];
              muxOutConnector[2] = fifoOut[4][12];
              muxOutConnector[3] = fifoOut[5][12];
              muxOutConnector[4] = fifoOut[6][12];
              muxOutConnector[5] = fifoOut[7][12];
              muxOutConnector[6] = fifoOut[8][12];
              muxOutConnector[7] = fifoOut[9][12];
              muxOutConnector[8] = fifoOut[10][12];
              muxOutConnector[9] = fifoOut[11][12];
              muxOutConnector[10] = fifoOut[12][12];
              muxOutConnector[11] = fifoOut[13][12];
              muxOutConnector[12] = fifoOut[14][12];
              muxOutConnector[13] = fifoOut[15][12];
              muxOutConnector[14] = fifoOut[16][12];
              muxOutConnector[15] = fifoOut[31][11];
              muxOutConnector[16] = fifoOut[32][11];
              muxOutConnector[17] = fifoOut[33][11];
              muxOutConnector[18] = fifoOut[34][11];
              muxOutConnector[19] = fifoOut[35][11];
              muxOutConnector[20] = fifoOut[36][11];
              muxOutConnector[21] = fifoOut[37][11];
              muxOutConnector[22] = fifoOut[38][11];
              muxOutConnector[23] = fifoOut[39][11];
              muxOutConnector[24] = fifoOut[40][11];
              muxOutConnector[25] = fifoOut[41][11];
              muxOutConnector[26] = fifoOut[3][8];
              muxOutConnector[27] = fifoOut[4][8];
              muxOutConnector[28] = fifoOut[5][8];
              muxOutConnector[29] = fifoOut[6][8];
              muxOutConnector[30] = fifoOut[7][8];
              muxOutConnector[31] = fifoOut[8][8];
              muxOutConnector[32] = fifoOut[9][8];
              muxOutConnector[33] = fifoOut[10][8];
              muxOutConnector[34] = fifoOut[11][8];
              muxOutConnector[35] = fifoOut[12][8];
              muxOutConnector[36] = fifoOut[13][8];
              muxOutConnector[37] = fifoOut[14][8];
              muxOutConnector[38] = fifoOut[15][8];
              muxOutConnector[39] = fifoOut[16][8];
              muxOutConnector[40] = fifoOut[17][8];
              muxOutConnector[41] = fifoOut[18][8];
              muxOutConnector[42] = fifoOut[19][8];
              muxOutConnector[43] = fifoOut[20][8];
              muxOutConnector[44] = fifoOut[21][8];
              muxOutConnector[45] = fifoOut[22][8];
              muxOutConnector[46] = fifoOut[23][8];
              muxOutConnector[47] = fifoOut[24][8];
              muxOutConnector[48] = fifoOut[25][8];
              muxOutConnector[49] = fifoOut[0][7];
              muxOutConnector[50] = fifoOut[1][7];
              muxOutConnector[51] = fifoOut[2][7];
       end
       13: begin
              muxOutConnector[0] = fifoOut[42][12];
              muxOutConnector[1] = fifoOut[43][12];
              muxOutConnector[2] = fifoOut[44][12];
              muxOutConnector[3] = fifoOut[45][12];
              muxOutConnector[4] = fifoOut[46][12];
              muxOutConnector[5] = fifoOut[47][12];
              muxOutConnector[6] = fifoOut[48][12];
              muxOutConnector[7] = fifoOut[49][12];
              muxOutConnector[8] = fifoOut[50][12];
              muxOutConnector[9] = fifoOut[51][12];
              muxOutConnector[10] = fifoOut[26][11];
              muxOutConnector[11] = fifoOut[27][11];
              muxOutConnector[12] = fifoOut[28][11];
              muxOutConnector[13] = fifoOut[29][11];
              muxOutConnector[14] = fifoOut[30][11];
              muxOutConnector[15] = fifoOut[31][11];
              muxOutConnector[16] = fifoOut[32][11];
              muxOutConnector[17] = fifoOut[33][11];
              muxOutConnector[18] = fifoOut[34][11];
              muxOutConnector[19] = fifoOut[35][11];
              muxOutConnector[20] = fifoOut[36][11];
              muxOutConnector[21] = fifoOut[37][11];
              muxOutConnector[22] = fifoOut[38][11];
              muxOutConnector[23] = fifoOut[39][11];
              muxOutConnector[24] = fifoOut[40][11];
              muxOutConnector[25] = fifoOut[41][11];
              muxOutConnector[26] = fifoOut[3][8];
              muxOutConnector[27] = fifoOut[4][8];
              muxOutConnector[28] = fifoOut[5][8];
              muxOutConnector[29] = fifoOut[6][8];
              muxOutConnector[30] = fifoOut[7][8];
              muxOutConnector[31] = fifoOut[8][8];
              muxOutConnector[32] = fifoOut[9][8];
              muxOutConnector[33] = fifoOut[10][8];
              muxOutConnector[34] = fifoOut[11][8];
              muxOutConnector[35] = fifoOut[12][8];
              muxOutConnector[36] = fifoOut[13][8];
              muxOutConnector[37] = fifoOut[14][8];
              muxOutConnector[38] = fifoOut[15][8];
              muxOutConnector[39] = fifoOut[16][8];
              muxOutConnector[40] = fifoOut[17][8];
              muxOutConnector[41] = fifoOut[18][8];
              muxOutConnector[42] = fifoOut[19][8];
              muxOutConnector[43] = fifoOut[20][8];
              muxOutConnector[44] = fifoOut[21][8];
              muxOutConnector[45] = fifoOut[22][8];
              muxOutConnector[46] = fifoOut[23][8];
              muxOutConnector[47] = fifoOut[24][8];
              muxOutConnector[48] = fifoOut[25][8];
              muxOutConnector[49] = fifoOut[0][7];
              muxOutConnector[50] = fifoOut[1][7];
              muxOutConnector[51] = fifoOut[2][7];
       end
       14: begin
              muxOutConnector[0] = fifoOut[42][12];
              muxOutConnector[1] = fifoOut[43][12];
              muxOutConnector[2] = fifoOut[44][12];
              muxOutConnector[3] = fifoOut[45][12];
              muxOutConnector[4] = fifoOut[46][12];
              muxOutConnector[5] = fifoOut[47][12];
              muxOutConnector[6] = fifoOut[48][12];
              muxOutConnector[7] = fifoOut[49][12];
              muxOutConnector[8] = fifoOut[50][12];
              muxOutConnector[9] = fifoOut[51][12];
              muxOutConnector[10] = fifoOut[26][11];
              muxOutConnector[11] = fifoOut[27][11];
              muxOutConnector[12] = fifoOut[28][11];
              muxOutConnector[13] = fifoOut[29][11];
              muxOutConnector[14] = fifoOut[30][11];
              muxOutConnector[15] = fifoOut[31][11];
              muxOutConnector[16] = fifoOut[32][11];
              muxOutConnector[17] = fifoOut[33][11];
              muxOutConnector[18] = fifoOut[34][11];
              muxOutConnector[19] = fifoOut[35][11];
              muxOutConnector[20] = fifoOut[36][11];
              muxOutConnector[21] = fifoOut[37][11];
              muxOutConnector[22] = fifoOut[38][11];
              muxOutConnector[23] = fifoOut[39][11];
              muxOutConnector[24] = fifoOut[40][11];
              muxOutConnector[25] = fifoOut[41][11];
              muxOutConnector[26] = fifoOut[3][8];
              muxOutConnector[27] = fifoOut[4][8];
              muxOutConnector[28] = fifoOut[5][8];
              muxOutConnector[29] = fifoOut[6][8];
              muxOutConnector[30] = fifoOut[7][8];
              muxOutConnector[31] = fifoOut[8][8];
              muxOutConnector[32] = fifoOut[9][8];
              muxOutConnector[33] = fifoOut[10][8];
              muxOutConnector[34] = fifoOut[11][8];
              muxOutConnector[35] = fifoOut[12][8];
              muxOutConnector[36] = fifoOut[13][8];
              muxOutConnector[37] = fifoOut[14][8];
              muxOutConnector[38] = fifoOut[15][8];
              muxOutConnector[39] = fifoOut[16][8];
              muxOutConnector[40] = fifoOut[17][8];
              muxOutConnector[41] = fifoOut[18][8];
              muxOutConnector[42] = fifoOut[19][8];
              muxOutConnector[43] = fifoOut[20][8];
              muxOutConnector[44] = fifoOut[21][8];
              muxOutConnector[45] = fifoOut[22][8];
              muxOutConnector[46] = fifoOut[23][8];
              muxOutConnector[47] = fifoOut[24][8];
              muxOutConnector[48] = fifoOut[25][8];
              muxOutConnector[49] = fifoOut[0][7];
              muxOutConnector[50] = fifoOut[1][7];
              muxOutConnector[51] = fifoOut[2][7];
       end
       15: begin
              muxOutConnector[0] = fifoOut[42][12];
              muxOutConnector[1] = fifoOut[43][12];
              muxOutConnector[2] = fifoOut[44][12];
              muxOutConnector[3] = fifoOut[45][12];
              muxOutConnector[4] = fifoOut[46][12];
              muxOutConnector[5] = fifoOut[47][12];
              muxOutConnector[6] = fifoOut[48][12];
              muxOutConnector[7] = fifoOut[49][12];
              muxOutConnector[8] = fifoOut[50][12];
              muxOutConnector[9] = fifoOut[51][12];
              muxOutConnector[10] = fifoOut[26][11];
              muxOutConnector[11] = fifoOut[27][11];
              muxOutConnector[12] = fifoOut[28][11];
              muxOutConnector[13] = fifoOut[29][11];
              muxOutConnector[14] = fifoOut[30][11];
              muxOutConnector[15] = fifoOut[31][11];
              muxOutConnector[16] = fifoOut[32][11];
              muxOutConnector[17] = fifoOut[33][11];
              muxOutConnector[18] = fifoOut[34][11];
              muxOutConnector[19] = fifoOut[35][11];
              muxOutConnector[20] = fifoOut[36][11];
              muxOutConnector[21] = fifoOut[37][11];
              muxOutConnector[22] = fifoOut[38][11];
              muxOutConnector[23] = fifoOut[39][11];
              muxOutConnector[24] = fifoOut[40][11];
              muxOutConnector[25] = fifoOut[41][11];
              muxOutConnector[26] = fifoOut[3][8];
              muxOutConnector[27] = fifoOut[4][8];
              muxOutConnector[28] = fifoOut[5][8];
              muxOutConnector[29] = fifoOut[6][8];
              muxOutConnector[30] = fifoOut[7][8];
              muxOutConnector[31] = fifoOut[8][8];
              muxOutConnector[32] = fifoOut[9][8];
              muxOutConnector[33] = fifoOut[10][8];
              muxOutConnector[34] = fifoOut[11][8];
              muxOutConnector[35] = fifoOut[12][8];
              muxOutConnector[36] = fifoOut[13][8];
              muxOutConnector[37] = fifoOut[14][8];
              muxOutConnector[38] = fifoOut[15][8];
              muxOutConnector[39] = fifoOut[16][8];
              muxOutConnector[40] = fifoOut[17][8];
              muxOutConnector[41] = fifoOut[18][8];
              muxOutConnector[42] = fifoOut[19][8];
              muxOutConnector[43] = fifoOut[20][8];
              muxOutConnector[44] = fifoOut[21][8];
              muxOutConnector[45] = fifoOut[22][8];
              muxOutConnector[46] = fifoOut[23][8];
              muxOutConnector[47] = fifoOut[24][8];
              muxOutConnector[48] = fifoOut[25][8];
              muxOutConnector[49] = fifoOut[0][7];
              muxOutConnector[50] = fifoOut[1][7];
              muxOutConnector[51] = fifoOut[2][7];
       end
       16: begin
              muxOutConnector[0] = fifoOut[42][12];
              muxOutConnector[1] = fifoOut[43][12];
              muxOutConnector[2] = fifoOut[44][12];
              muxOutConnector[3] = fifoOut[45][12];
              muxOutConnector[4] = fifoOut[46][12];
              muxOutConnector[5] = fifoOut[47][12];
              muxOutConnector[6] = fifoOut[48][12];
              muxOutConnector[7] = fifoOut[49][12];
              muxOutConnector[8] = fifoOut[50][12];
              muxOutConnector[9] = fifoOut[51][12];
              muxOutConnector[10] = fifoOut[26][11];
              muxOutConnector[11] = fifoOut[27][11];
              muxOutConnector[12] = fifoOut[28][11];
              muxOutConnector[13] = fifoOut[29][11];
              muxOutConnector[14] = fifoOut[30][11];
              muxOutConnector[15] = fifoOut[31][11];
              muxOutConnector[16] = fifoOut[32][11];
              muxOutConnector[17] = fifoOut[33][11];
              muxOutConnector[18] = fifoOut[34][11];
              muxOutConnector[19] = fifoOut[35][11];
              muxOutConnector[20] = fifoOut[36][11];
              muxOutConnector[21] = fifoOut[37][11];
              muxOutConnector[22] = fifoOut[38][11];
              muxOutConnector[23] = fifoOut[39][11];
              muxOutConnector[24] = fifoOut[40][11];
              muxOutConnector[25] = fifoOut[41][11];
              muxOutConnector[26] = fifoOut[3][8];
              muxOutConnector[27] = fifoOut[4][8];
              muxOutConnector[28] = fifoOut[5][8];
              muxOutConnector[29] = fifoOut[6][8];
              muxOutConnector[30] = fifoOut[7][8];
              muxOutConnector[31] = fifoOut[8][8];
              muxOutConnector[32] = fifoOut[9][8];
              muxOutConnector[33] = fifoOut[10][8];
              muxOutConnector[34] = fifoOut[11][8];
              muxOutConnector[35] = fifoOut[12][8];
              muxOutConnector[36] = fifoOut[13][8];
              muxOutConnector[37] = fifoOut[14][8];
              muxOutConnector[38] = fifoOut[15][8];
              muxOutConnector[39] = fifoOut[16][8];
              muxOutConnector[40] = fifoOut[17][8];
              muxOutConnector[41] = fifoOut[18][8];
              muxOutConnector[42] = fifoOut[19][8];
              muxOutConnector[43] = fifoOut[20][8];
              muxOutConnector[44] = fifoOut[21][8];
              muxOutConnector[45] = fifoOut[22][8];
              muxOutConnector[46] = fifoOut[23][8];
              muxOutConnector[47] = fifoOut[24][8];
              muxOutConnector[48] = fifoOut[25][8];
              muxOutConnector[49] = fifoOut[0][7];
              muxOutConnector[50] = fifoOut[1][7];
              muxOutConnector[51] = fifoOut[2][7];
       end
       17: begin
              muxOutConnector[0] = fifoOut[42][12];
              muxOutConnector[1] = fifoOut[43][12];
              muxOutConnector[2] = fifoOut[44][12];
              muxOutConnector[3] = fifoOut[45][12];
              muxOutConnector[4] = fifoOut[46][12];
              muxOutConnector[5] = fifoOut[47][12];
              muxOutConnector[6] = fifoOut[48][12];
              muxOutConnector[7] = fifoOut[49][12];
              muxOutConnector[8] = fifoOut[50][12];
              muxOutConnector[9] = fifoOut[51][12];
              muxOutConnector[10] = fifoOut[26][11];
              muxOutConnector[11] = fifoOut[27][11];
              muxOutConnector[12] = fifoOut[28][11];
              muxOutConnector[13] = fifoOut[29][11];
              muxOutConnector[14] = fifoOut[30][11];
              muxOutConnector[15] = fifoOut[31][11];
              muxOutConnector[16] = fifoOut[32][11];
              muxOutConnector[17] = fifoOut[33][11];
              muxOutConnector[18] = fifoOut[34][11];
              muxOutConnector[19] = fifoOut[35][11];
              muxOutConnector[20] = fifoOut[36][11];
              muxOutConnector[21] = fifoOut[37][11];
              muxOutConnector[22] = fifoOut[38][11];
              muxOutConnector[23] = fifoOut[39][11];
              muxOutConnector[24] = fifoOut[40][11];
              muxOutConnector[25] = fifoOut[41][11];
              muxOutConnector[26] = fifoOut[3][8];
              muxOutConnector[27] = fifoOut[4][8];
              muxOutConnector[28] = fifoOut[5][8];
              muxOutConnector[29] = fifoOut[6][8];
              muxOutConnector[30] = fifoOut[7][8];
              muxOutConnector[31] = fifoOut[8][8];
              muxOutConnector[32] = fifoOut[9][8];
              muxOutConnector[33] = fifoOut[10][8];
              muxOutConnector[34] = fifoOut[11][8];
              muxOutConnector[35] = fifoOut[12][8];
              muxOutConnector[36] = fifoOut[13][8];
              muxOutConnector[37] = fifoOut[14][8];
              muxOutConnector[38] = fifoOut[15][8];
              muxOutConnector[39] = fifoOut[16][8];
              muxOutConnector[40] = fifoOut[17][8];
              muxOutConnector[41] = fifoOut[18][8];
              muxOutConnector[42] = fifoOut[19][8];
              muxOutConnector[43] = fifoOut[20][8];
              muxOutConnector[44] = fifoOut[21][8];
              muxOutConnector[45] = fifoOut[22][8];
              muxOutConnector[46] = fifoOut[23][8];
              muxOutConnector[47] = fifoOut[24][8];
              muxOutConnector[48] = fifoOut[25][8];
              muxOutConnector[49] = fifoOut[0][7];
              muxOutConnector[50] = fifoOut[1][7];
              muxOutConnector[51] = fifoOut[2][7];
       end
       18: begin
              muxOutConnector[0] = fifoOut[42][12];
              muxOutConnector[1] = fifoOut[43][12];
              muxOutConnector[2] = fifoOut[44][12];
              muxOutConnector[3] = fifoOut[45][12];
              muxOutConnector[4] = fifoOut[46][12];
              muxOutConnector[5] = fifoOut[47][12];
              muxOutConnector[6] = fifoOut[48][12];
              muxOutConnector[7] = fifoOut[49][12];
              muxOutConnector[8] = fifoOut[50][12];
              muxOutConnector[9] = fifoOut[51][12];
              muxOutConnector[10] = fifoOut[26][11];
              muxOutConnector[11] = fifoOut[27][11];
              muxOutConnector[12] = fifoOut[28][11];
              muxOutConnector[13] = fifoOut[29][11];
              muxOutConnector[14] = fifoOut[30][11];
              muxOutConnector[15] = fifoOut[31][11];
              muxOutConnector[16] = fifoOut[32][11];
              muxOutConnector[17] = fifoOut[33][11];
              muxOutConnector[18] = fifoOut[34][11];
              muxOutConnector[19] = fifoOut[35][11];
              muxOutConnector[20] = fifoOut[36][11];
              muxOutConnector[21] = fifoOut[37][11];
              muxOutConnector[22] = fifoOut[38][11];
              muxOutConnector[23] = fifoOut[39][11];
              muxOutConnector[24] = fifoOut[40][11];
              muxOutConnector[25] = fifoOut[41][11];
              muxOutConnector[26] = fifoOut[3][8];
              muxOutConnector[27] = fifoOut[4][8];
              muxOutConnector[28] = fifoOut[5][8];
              muxOutConnector[29] = fifoOut[6][8];
              muxOutConnector[30] = fifoOut[7][8];
              muxOutConnector[31] = fifoOut[8][8];
              muxOutConnector[32] = fifoOut[9][8];
              muxOutConnector[33] = fifoOut[10][8];
              muxOutConnector[34] = fifoOut[11][8];
              muxOutConnector[35] = fifoOut[12][8];
              muxOutConnector[36] = fifoOut[13][8];
              muxOutConnector[37] = fifoOut[14][8];
              muxOutConnector[38] = fifoOut[15][8];
              muxOutConnector[39] = fifoOut[16][8];
              muxOutConnector[40] = fifoOut[17][8];
              muxOutConnector[41] = fifoOut[18][8];
              muxOutConnector[42] = fifoOut[19][8];
              muxOutConnector[43] = fifoOut[20][8];
              muxOutConnector[44] = fifoOut[21][8];
              muxOutConnector[45] = fifoOut[22][8];
              muxOutConnector[46] = fifoOut[23][8];
              muxOutConnector[47] = fifoOut[24][8];
              muxOutConnector[48] = fifoOut[25][8];
              muxOutConnector[49] = fifoOut[0][7];
              muxOutConnector[50] = fifoOut[1][7];
              muxOutConnector[51] = fifoOut[2][7];
       end
       19: begin
              muxOutConnector[0] = fifoOut[42][12];
              muxOutConnector[1] = fifoOut[43][12];
              muxOutConnector[2] = fifoOut[44][12];
              muxOutConnector[3] = fifoOut[45][12];
              muxOutConnector[4] = fifoOut[46][12];
              muxOutConnector[5] = fifoOut[47][12];
              muxOutConnector[6] = fifoOut[48][12];
              muxOutConnector[7] = fifoOut[49][12];
              muxOutConnector[8] = fifoOut[50][12];
              muxOutConnector[9] = fifoOut[51][12];
              muxOutConnector[10] = fifoOut[26][11];
              muxOutConnector[11] = fifoOut[27][11];
              muxOutConnector[12] = fifoOut[28][11];
              muxOutConnector[13] = fifoOut[29][11];
              muxOutConnector[14] = fifoOut[30][11];
              muxOutConnector[15] = fifoOut[31][11];
              muxOutConnector[16] = fifoOut[32][11];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[3][8];
              muxOutConnector[27] = fifoOut[4][8];
              muxOutConnector[28] = fifoOut[5][8];
              muxOutConnector[29] = fifoOut[6][8];
              muxOutConnector[30] = fifoOut[7][8];
              muxOutConnector[31] = fifoOut[8][8];
              muxOutConnector[32] = fifoOut[9][8];
              muxOutConnector[33] = fifoOut[10][8];
              muxOutConnector[34] = fifoOut[11][8];
              muxOutConnector[35] = fifoOut[12][8];
              muxOutConnector[36] = fifoOut[13][8];
              muxOutConnector[37] = fifoOut[14][8];
              muxOutConnector[38] = fifoOut[15][8];
              muxOutConnector[39] = fifoOut[16][8];
              muxOutConnector[40] = fifoOut[17][8];
              muxOutConnector[41] = fifoOut[18][8];
              muxOutConnector[42] = fifoOut[19][8];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
