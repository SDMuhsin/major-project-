`timescale 1ns / 1ps
module Dmem_circ2_scripted(
		 muxOut,
		 dMemIn,
		 wr_en,
		 reaccessAddress,
		 reaccess_lyr,
		 rd_en, clk, rst 
 );
parameter r = 52;
parameter c = 12;
parameter w = 6;
parameter ADDRESSWIDTH = 5;

parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 
output wire [r*w -1 : 0]muxOut;// r numbers of w bits
input [r*w-1:0]dMemIn;
input wr_en;
input [ADDRESSWIDTH-1:0]reaccessAddress;
input reaccess_lyr;
input rd_en;
input clk,rst;

wire [(ADDRESSWIDTH+1)-1:0]case_sel;//{layer,address}
wire [w-1:0]dMemInDummy[r-1:0];
reg [w-1:0]muxOutWire[r-1:0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<r;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutWire[k];
        assign dMemInDummy[k] = dMemIn[ (k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always @(posedge clk) begin
    if (rst) begin
         for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] = 0;
           end
        end
    end
    else begin
    if(wr_en) begin
        // Set (i,j)th value = (i,j-1)th value
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Load Inputs
        for(i = r-1; i > -1; i=i-1) begin
            fifoOut[i][0] <= dMemInDummy[i]; 
        end
    end
    else begin 
        // Set (i,j)th value = (i,j)th value
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <= fifoOut[i][j];
            end
        end
    end
    end
end

assign case_sel = rd_en ? {reaccess_lyr,reaccessAddress} : {1'd1,READDISABLEDCASE};

always@(*) begin
    case(case_sel)

		 {1'd0, 5'd0} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd1} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd2} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd3} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd4} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd5} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd6} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = fifoOut[ 0 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 1 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 2 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 3 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 4 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 5 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 6 ][ 3 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 7 ][ 3 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 8 ][ 3 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 9 ][ 3 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 10 ][ 3 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 11 ][ 3 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 12 ][ 3 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 13 ][ 3 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 14 ][ 3 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 15 ][ 3 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 16 ][ 3 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 22 ][ 3 ]; 
		 end
		 {1'd0, 5'd7} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 23 ][ 4 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 24 ][ 4 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 25 ][ 4 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 0 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 1 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 2 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 3 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 4 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 5 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 6 ][ 3 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 7 ][ 3 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 8 ][ 3 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 9 ][ 3 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 10 ][ 3 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 11 ][ 3 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 12 ][ 3 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 13 ][ 3 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 14 ][ 3 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 15 ][ 3 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 16 ][ 3 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 22 ][ 3 ]; 
		 end
		 {1'd0, 5'd8} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 23 ][ 4 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 24 ][ 4 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 25 ][ 4 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 0 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 1 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 2 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 3 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 4 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 5 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 6 ][ 3 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 7 ][ 3 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 8 ][ 3 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 9 ][ 3 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 10 ][ 3 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 11 ][ 3 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 12 ][ 3 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 13 ][ 3 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 14 ][ 3 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 15 ][ 3 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 16 ][ 3 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 22 ][ 3 ]; 
		 end
		 {1'd0, 5'd9} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 23 ][ 4 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 24 ][ 4 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 25 ][ 4 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 0 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 1 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 2 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 3 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 4 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 5 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 6 ][ 3 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 7 ][ 3 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 8 ][ 3 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 9 ][ 3 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 10 ][ 3 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 11 ][ 3 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 12 ][ 3 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 13 ][ 3 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 14 ][ 3 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 15 ][ 3 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 16 ][ 3 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 22 ][ 3 ]; 
		 end
		 {1'd0, 5'd10} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 23 ][ 4 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 24 ][ 4 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 25 ][ 4 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 0 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 1 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 2 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 3 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 4 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 5 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 6 ][ 3 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 7 ][ 3 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 8 ][ 3 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 9 ][ 3 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 10 ][ 3 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 11 ][ 3 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 12 ][ 3 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 13 ][ 3 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 14 ][ 3 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 15 ][ 3 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 16 ][ 3 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 22 ][ 3 ]; 
		 end
		 {1'd0, 5'd11} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 23 ][ 4 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 24 ][ 4 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 25 ][ 4 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 0 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 1 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 2 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 3 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 4 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 5 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 6 ][ 3 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 7 ][ 3 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 8 ][ 3 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 9 ][ 3 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 10 ][ 3 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 11 ][ 3 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 12 ][ 3 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 13 ][ 3 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 14 ][ 3 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 15 ][ 3 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 16 ][ 3 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 22 ][ 3 ]; 
		 end
		 {1'd0, 5'd12} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 23 ][ 4 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 24 ][ 4 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 25 ][ 4 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 0 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 1 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 2 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 3 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 4 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 5 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 6 ][ 3 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 7 ][ 3 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 8 ][ 3 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 9 ][ 3 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 10 ][ 3 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 11 ][ 3 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 12 ][ 3 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 13 ][ 3 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 14 ][ 3 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 15 ][ 3 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 16 ][ 3 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 22 ][ 3 ]; 
		 end
		 {1'd0, 5'd13} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = fifoOut[ 26 ][ 10 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 27 ][ 10 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 28 ][ 10 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 29 ][ 10 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 30 ][ 10 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 31 ][ 10 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 32 ][ 10 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 33 ][ 10 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 34 ][ 10 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 35 ][ 10 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 36 ][ 10 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 37 ][ 10 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 23 ][ 4 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 24 ][ 4 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 25 ][ 4 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 0 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 1 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 2 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 3 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 4 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 5 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 6 ][ 3 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 7 ][ 3 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 8 ][ 3 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 9 ][ 3 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 10 ][ 3 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 11 ][ 3 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 12 ][ 3 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 13 ][ 3 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 14 ][ 3 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 15 ][ 3 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 16 ][ 3 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 22 ][ 3 ]; 
		 end
		 {1'd0, 5'd14} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 38 ][ 11 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 39 ][ 11 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 40 ][ 11 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 41 ][ 11 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 42 ][ 11 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 43 ][ 11 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 44 ][ 11 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 45 ][ 11 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 46 ][ 11 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 47 ][ 11 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 48 ][ 11 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 49 ][ 11 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 50 ][ 11 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 51 ][ 11 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 26 ][ 10 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 27 ][ 10 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 28 ][ 10 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 29 ][ 10 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 30 ][ 10 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 31 ][ 10 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 32 ][ 10 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 33 ][ 10 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 34 ][ 10 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 35 ][ 10 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 36 ][ 10 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 37 ][ 10 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 23 ][ 4 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 24 ][ 4 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 25 ][ 4 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 0 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 1 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 2 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 3 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 4 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 5 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 6 ][ 3 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 7 ][ 3 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 8 ][ 3 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 9 ][ 3 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 10 ][ 3 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 11 ][ 3 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 12 ][ 3 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 13 ][ 3 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 14 ][ 3 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 15 ][ 3 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 16 ][ 3 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 22 ][ 3 ]; 
		 end
		 {1'd0, 5'd15} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 38 ][ 11 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 39 ][ 11 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 40 ][ 11 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 41 ][ 11 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 42 ][ 11 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 43 ][ 11 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 44 ][ 11 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 45 ][ 11 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 46 ][ 11 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 47 ][ 11 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 48 ][ 11 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 49 ][ 11 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 50 ][ 11 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 51 ][ 11 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 26 ][ 10 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 27 ][ 10 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 28 ][ 10 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 29 ][ 10 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 30 ][ 10 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 31 ][ 10 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 32 ][ 10 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 33 ][ 10 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 34 ][ 10 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 35 ][ 10 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 36 ][ 10 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 37 ][ 10 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 23 ][ 4 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 24 ][ 4 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 25 ][ 4 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 0 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 1 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 2 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 3 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 4 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 5 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 6 ][ 3 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 7 ][ 3 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 8 ][ 3 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 9 ][ 3 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 10 ][ 3 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 11 ][ 3 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 12 ][ 3 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 13 ][ 3 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 14 ][ 3 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 15 ][ 3 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 16 ][ 3 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 22 ][ 3 ]; 
		 end
		 {1'd0, 5'd16} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 38 ][ 11 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 39 ][ 11 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 40 ][ 11 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 41 ][ 11 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 42 ][ 11 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 43 ][ 11 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 44 ][ 11 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 45 ][ 11 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 46 ][ 11 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 47 ][ 11 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 48 ][ 11 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 49 ][ 11 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 50 ][ 11 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 51 ][ 11 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 26 ][ 10 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 27 ][ 10 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 28 ][ 10 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 29 ][ 10 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 30 ][ 10 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 31 ][ 10 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 32 ][ 10 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 33 ][ 10 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 34 ][ 10 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 35 ][ 10 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 36 ][ 10 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 37 ][ 10 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 23 ][ 4 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 24 ][ 4 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 25 ][ 4 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 0 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 1 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 2 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 3 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 4 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 5 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 6 ][ 3 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 7 ][ 3 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 8 ][ 3 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 9 ][ 3 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 10 ][ 3 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 11 ][ 3 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 12 ][ 3 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 13 ][ 3 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 14 ][ 3 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 15 ][ 3 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 16 ][ 3 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 22 ][ 3 ]; 
		 end
		 {1'd0, 5'd17} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 38 ][ 11 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 39 ][ 11 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 40 ][ 11 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 41 ][ 11 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 42 ][ 11 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 43 ][ 11 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 44 ][ 11 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 45 ][ 11 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 46 ][ 11 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 47 ][ 11 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 48 ][ 11 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 49 ][ 11 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 50 ][ 11 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 51 ][ 11 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 26 ][ 10 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 27 ][ 10 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 28 ][ 10 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 29 ][ 10 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 30 ][ 10 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 31 ][ 10 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 32 ][ 10 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 33 ][ 10 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 34 ][ 10 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 35 ][ 10 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 36 ][ 10 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 37 ][ 10 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 23 ][ 4 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 24 ][ 4 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 25 ][ 4 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 0 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 1 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 2 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 3 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 4 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 5 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 6 ][ 3 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 7 ][ 3 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 8 ][ 3 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 9 ][ 3 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 10 ][ 3 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 11 ][ 3 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 12 ][ 3 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 13 ][ 3 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 14 ][ 3 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 15 ][ 3 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 16 ][ 3 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 22 ][ 3 ]; 
		 end
		 {1'd0, 5'd18} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 38 ][ 11 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 39 ][ 11 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 40 ][ 11 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 41 ][ 11 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 42 ][ 11 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 43 ][ 11 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 44 ][ 11 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 45 ][ 11 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 46 ][ 11 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 47 ][ 11 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 48 ][ 11 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 49 ][ 11 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 50 ][ 11 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 51 ][ 11 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 26 ][ 10 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 27 ][ 10 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 28 ][ 10 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 29 ][ 10 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 30 ][ 10 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 31 ][ 10 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 32 ][ 10 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 33 ][ 10 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 34 ][ 10 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 35 ][ 10 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 36 ][ 10 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 37 ][ 10 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 23 ][ 4 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 24 ][ 4 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 25 ][ 4 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 0 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 1 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 2 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 3 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 4 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 5 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 6 ][ 3 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 7 ][ 3 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 8 ][ 3 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 9 ][ 3 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 10 ][ 3 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 11 ][ 3 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 12 ][ 3 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 13 ][ 3 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 14 ][ 3 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 15 ][ 3 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 16 ][ 3 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 17 ][ 3 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 18 ][ 3 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 19 ][ 3 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 20 ][ 3 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 21 ][ 3 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 22 ][ 3 ]; 
		 end
		 {1'd0, 5'd19} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 38 ][ 11 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 39 ][ 11 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 40 ][ 11 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 41 ][ 11 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 42 ][ 11 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 43 ][ 11 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 44 ][ 11 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 45 ][ 11 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 46 ][ 11 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 47 ][ 11 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 48 ][ 11 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 49 ][ 11 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 50 ][ 11 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 51 ][ 11 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 26 ][ 10 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 27 ][ 10 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 28 ][ 10 ]; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 23 ][ 4 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 24 ][ 4 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 25 ][ 4 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 0 ][ 3 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 1 ][ 3 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 2 ][ 3 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 3 ][ 3 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 4 ][ 3 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 5 ][ 3 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 6 ][ 3 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 7 ][ 3 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 8 ][ 3 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 9 ][ 3 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 10 ][ 3 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 11 ][ 3 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 12 ][ 3 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 13 ][ 3 ]; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd0} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd1} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd2} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd3} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd4} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd5} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd6} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd7} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd8} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd9} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 31 ][ 6 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 32 ][ 6 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 33 ][ 6 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 34 ][ 6 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 35 ][ 6 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 36 ][ 6 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 37 ][ 6 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 38 ][ 6 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 39 ][ 6 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 40 ][ 6 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 41 ][ 6 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 42 ][ 6 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 43 ][ 6 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 44 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 45 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 46 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 47 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 48 ][ 6 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd10} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 31 ][ 6 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 32 ][ 6 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 33 ][ 6 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 34 ][ 6 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 35 ][ 6 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 36 ][ 6 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 37 ][ 6 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 38 ][ 6 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 39 ][ 6 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 40 ][ 6 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 41 ][ 6 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 42 ][ 6 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 43 ][ 6 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 44 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 45 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 46 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 47 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 48 ][ 6 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = fifoOut[ 0 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 1 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 2 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 3 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 11 ][ 7 ]; 
		 end
		 {1'd1, 5'd11} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 31 ][ 6 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 32 ][ 6 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 33 ][ 6 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 34 ][ 6 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 35 ][ 6 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 36 ][ 6 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 37 ][ 6 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 38 ][ 6 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 39 ][ 6 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 40 ][ 6 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 41 ][ 6 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 42 ][ 6 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 43 ][ 6 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 44 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 45 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 46 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 47 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 48 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 12 ][ 8 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 13 ][ 8 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 14 ][ 8 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 15 ][ 8 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 16 ][ 8 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 17 ][ 8 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 18 ][ 8 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 19 ][ 8 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 20 ][ 8 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 21 ][ 8 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 22 ][ 8 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 23 ][ 8 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 24 ][ 8 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 25 ][ 8 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 0 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 1 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 2 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 3 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 11 ][ 7 ]; 
		 end
		 {1'd1, 5'd12} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 31 ][ 6 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 32 ][ 6 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 33 ][ 6 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 34 ][ 6 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 35 ][ 6 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 36 ][ 6 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 37 ][ 6 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 38 ][ 6 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 39 ][ 6 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 40 ][ 6 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 41 ][ 6 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 42 ][ 6 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 43 ][ 6 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 44 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 45 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 46 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 47 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 48 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 12 ][ 8 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 13 ][ 8 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 14 ][ 8 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 15 ][ 8 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 16 ][ 8 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 17 ][ 8 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 18 ][ 8 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 19 ][ 8 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 20 ][ 8 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 21 ][ 8 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 22 ][ 8 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 23 ][ 8 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 24 ][ 8 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 25 ][ 8 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 0 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 1 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 2 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 3 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 11 ][ 7 ]; 
		 end
		 {1'd1, 5'd13} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 31 ][ 6 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 32 ][ 6 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 33 ][ 6 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 34 ][ 6 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 35 ][ 6 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 36 ][ 6 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 37 ][ 6 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 38 ][ 6 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 39 ][ 6 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 40 ][ 6 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 41 ][ 6 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 42 ][ 6 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 43 ][ 6 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 44 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 45 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 46 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 47 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 48 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 12 ][ 8 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 13 ][ 8 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 14 ][ 8 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 15 ][ 8 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 16 ][ 8 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 17 ][ 8 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 18 ][ 8 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 19 ][ 8 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 20 ][ 8 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 21 ][ 8 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 22 ][ 8 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 23 ][ 8 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 24 ][ 8 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 25 ][ 8 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 0 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 1 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 2 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 3 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 11 ][ 7 ]; 
		 end
		 {1'd1, 5'd14} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 31 ][ 6 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 32 ][ 6 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 33 ][ 6 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 34 ][ 6 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 35 ][ 6 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 36 ][ 6 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 37 ][ 6 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 38 ][ 6 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 39 ][ 6 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 40 ][ 6 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 41 ][ 6 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 42 ][ 6 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 43 ][ 6 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 44 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 45 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 46 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 47 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 48 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 12 ][ 8 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 13 ][ 8 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 14 ][ 8 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 15 ][ 8 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 16 ][ 8 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 17 ][ 8 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 18 ][ 8 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 19 ][ 8 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 20 ][ 8 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 21 ][ 8 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 22 ][ 8 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 23 ][ 8 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 24 ][ 8 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 25 ][ 8 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 0 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 1 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 2 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 3 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 11 ][ 7 ]; 
		 end
		 {1'd1, 5'd15} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 31 ][ 6 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 32 ][ 6 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 33 ][ 6 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 34 ][ 6 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 35 ][ 6 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 36 ][ 6 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 37 ][ 6 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 38 ][ 6 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 39 ][ 6 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 40 ][ 6 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 41 ][ 6 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 42 ][ 6 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 43 ][ 6 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 44 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 45 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 46 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 47 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 48 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 12 ][ 8 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 13 ][ 8 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 14 ][ 8 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 15 ][ 8 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 16 ][ 8 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 17 ][ 8 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 18 ][ 8 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 19 ][ 8 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 20 ][ 8 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 21 ][ 8 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 22 ][ 8 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 23 ][ 8 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 24 ][ 8 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 25 ][ 8 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 0 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 1 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 2 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 3 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 11 ][ 7 ]; 
		 end
		 {1'd1, 5'd16} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 31 ][ 6 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 32 ][ 6 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 33 ][ 6 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 34 ][ 6 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 35 ][ 6 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 36 ][ 6 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 37 ][ 6 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 38 ][ 6 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 39 ][ 6 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 40 ][ 6 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 41 ][ 6 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 42 ][ 6 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 43 ][ 6 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 44 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 45 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 46 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 47 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 48 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 12 ][ 8 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 13 ][ 8 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 14 ][ 8 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 15 ][ 8 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 16 ][ 8 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 17 ][ 8 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 18 ][ 8 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 19 ][ 8 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 20 ][ 8 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 21 ][ 8 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 22 ][ 8 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 23 ][ 8 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 24 ][ 8 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 25 ][ 8 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 0 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 1 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 2 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 3 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 11 ][ 7 ]; 
		 end
		 {1'd1, 5'd17} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 31 ][ 6 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 32 ][ 6 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 33 ][ 6 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 34 ][ 6 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 35 ][ 6 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 36 ][ 6 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 37 ][ 6 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 38 ][ 6 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 39 ][ 6 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 40 ][ 6 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 41 ][ 6 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 42 ][ 6 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 43 ][ 6 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 44 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 45 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 46 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 47 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 48 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 12 ][ 8 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 13 ][ 8 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 14 ][ 8 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 15 ][ 8 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 16 ][ 8 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 17 ][ 8 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 18 ][ 8 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 19 ][ 8 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 20 ][ 8 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 21 ][ 8 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 22 ][ 8 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 23 ][ 8 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 24 ][ 8 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 25 ][ 8 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 0 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 1 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 2 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 3 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 11 ][ 7 ]; 
		 end
		 {1'd1, 5'd18} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 31 ][ 6 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 32 ][ 6 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 33 ][ 6 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 34 ][ 6 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 35 ][ 6 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 36 ][ 6 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 37 ][ 6 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 38 ][ 6 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 39 ][ 6 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 40 ][ 6 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 41 ][ 6 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 42 ][ 6 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 43 ][ 6 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 44 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 45 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 46 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 47 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 48 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 12 ][ 8 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 13 ][ 8 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 14 ][ 8 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 15 ][ 8 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 16 ][ 8 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 17 ][ 8 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 18 ][ 8 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 19 ][ 8 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 20 ][ 8 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 21 ][ 8 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 22 ][ 8 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 23 ][ 8 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 24 ][ 8 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 25 ][ 8 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 0 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 1 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 2 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 3 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 11 ][ 7 ]; 
		 end
		 {1'd1, 5'd19} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 31 ][ 6 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 32 ][ 6 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 33 ][ 6 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 34 ][ 6 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 35 ][ 6 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 36 ][ 6 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 37 ][ 6 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 38 ][ 6 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 39 ][ 6 ]; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 12 ][ 8 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 13 ][ 8 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 14 ][ 8 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 15 ][ 8 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 16 ][ 8 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 17 ][ 8 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 18 ][ 8 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 19 ][ 8 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 20 ][ 8 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 21 ][ 8 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 22 ][ 8 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 23 ][ 8 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 24 ][ 8 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 25 ][ 8 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 0 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 1 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 2 ][ 7 ]; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
    default:begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
    end
    endcase
end
endmodule
