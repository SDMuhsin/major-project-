`timescale 1ns / 1ps
module Dmem_circ13_scripted(
		 muxOut,
		 dMemIn,
		 wr_en,
		 reaccessAddress,
		 reaccess_lyr,
		 rd_en, clk, rst 
 );
parameter r = 52;
parameter c = 14;
parameter w = 6;
parameter ADDRESSWIDTH = 5;

parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 
output wire [r*w -1 : 0]muxOut;// r numbers of w bits
input [r*w-1:0]dMemIn;
input wr_en;
input [ADDRESSWIDTH-1:0]reaccessAddress;
input reaccess_lyr;
input rd_en;
input clk,rst;

wire [(ADDRESSWIDTH+1)-1:0]case_sel;//{layer,address}
wire [w-1:0]dMemInDummy[r-1:0];
reg [w-1:0]muxOutWire[r-1:0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<r;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutWire[k];
        assign dMemInDummy[k] = dMemIn[ (k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always @(posedge clk) begin
    if (!rst) begin
         for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] = 0;
           end
        end
    end
    else begin
    if(wr_en) begin
        // Set (i,j)th value = (i,j-1)th value
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Load Inputs
        for(i = r-1; i > -1; i=i-1) begin
            fifoOut[i][0] <= dMemInDummy[i]; 
        end
    end
    else begin 
        // Set (i,j)th value = (i,j)th value
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <= fifoOut[i][j];
            end
        end
    end
    end
end

assign case_sel = rd_en ? {reaccess_lyr,reaccessAddress} : {1'd1,READDISABLEDCASE};

always@(*) begin
    case(case_sel)

		 {1'd0, 5'd0} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd1} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd2} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd3} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd4} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd5} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd6} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd7} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd8} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd0, 5'd9} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 6 ]; 
		 end
		 {1'd0, 5'd10} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 7 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 7 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 7 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 7 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 7 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 7 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 7 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 7 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 7 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 7 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 7 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 7 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 7 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 7 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 7 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 7 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 7 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 7 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 6 ]; 
		 end
		 {1'd0, 5'd11} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 7 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 7 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 7 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 7 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 7 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 7 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 7 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 7 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 7 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 7 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 7 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 7 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 7 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 7 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 7 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 7 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 7 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 7 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 6 ]; 
		 end
		 {1'd0, 5'd12} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 7 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 7 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 7 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 7 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 7 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 7 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 7 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 7 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 7 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 7 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 7 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 7 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 7 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 7 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 7 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 7 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 7 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 7 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 6 ]; 
		 end
		 {1'd0, 5'd13} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 7 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 7 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 7 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 7 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 7 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 7 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 7 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 7 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 7 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 7 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 7 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 7 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 7 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 7 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 7 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 7 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 7 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 7 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 6 ]; 
		 end
		 {1'd0, 5'd14} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 7 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 7 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 7 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 7 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 7 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 7 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 7 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 7 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 7 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 7 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 7 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 7 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 7 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 7 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 7 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 7 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 7 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 7 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 6 ]; 
		 end
		 {1'd0, 5'd15} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 7 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 7 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 7 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 7 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 7 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 7 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 7 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 7 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 7 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 7 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 7 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 7 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 7 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 7 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 7 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 7 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 7 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 7 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 6 ]; 
		 end
		 {1'd0, 5'd16} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 7 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 7 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 7 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 7 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 7 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 7 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 7 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 7 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 7 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 7 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 7 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 7 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 7 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 7 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 7 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 7 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 7 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 7 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 6 ]; 
		 end
		 {1'd0, 5'd17} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 7 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 7 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 7 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 7 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 7 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 7 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 7 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 7 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 7 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 7 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 7 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 7 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 7 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 7 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 7 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 7 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 7 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 7 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 6 ]; 
		 end
		 {1'd0, 5'd18} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 7 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 7 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 7 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 7 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 7 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 7 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 7 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 7 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 7 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 7 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 7 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 7 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 48 ][ 7 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 49 ][ 7 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 50 ][ 7 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 51 ][ 7 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 26 ][ 6 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 27 ][ 6 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 28 ][ 6 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 29 ][ 6 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 30 ][ 6 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 7 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 7 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 7 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 7 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 7 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 7 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 7 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 7 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 21 ][ 7 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 22 ][ 7 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 23 ][ 7 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 24 ][ 7 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 25 ][ 7 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 0 ][ 6 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 1 ][ 6 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 2 ][ 6 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 3 ][ 6 ]; 
		 end
		 {1'd0, 5'd19} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 31 ][ 7 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 32 ][ 7 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 33 ][ 7 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 34 ][ 7 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 35 ][ 7 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 36 ][ 7 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 37 ][ 7 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 38 ][ 7 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 39 ][ 7 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 40 ][ 7 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 41 ][ 7 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 42 ][ 7 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 43 ][ 7 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 44 ][ 7 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 45 ][ 7 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 46 ][ 7 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 47 ][ 7 ]; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 4 ][ 7 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 5 ][ 7 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 6 ][ 7 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 7 ][ 7 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 8 ][ 7 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 9 ][ 7 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 10 ][ 7 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 11 ][ 7 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 12 ][ 7 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 13 ][ 7 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 14 ][ 7 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 15 ][ 7 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 16 ][ 7 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 17 ][ 7 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 18 ][ 7 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 19 ][ 7 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 20 ][ 7 ]; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd0} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd1} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd2} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd3} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd4} : begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd5} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd6} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd7} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd8} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd9} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd10} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd11} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd12} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd13} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd14} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
		 {1'd1, 5'd15} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = fifoOut[ 0 ][ 12 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 1 ][ 12 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 2 ][ 12 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 3 ][ 12 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 4 ][ 12 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 5 ][ 12 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 6 ][ 12 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 7 ][ 12 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 8 ][ 12 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 9 ][ 12 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 10 ][ 12 ]; 
		 end
		 {1'd1, 5'd16} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 11 ][ 13 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 12 ][ 13 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 13 ][ 13 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 14 ][ 13 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 15 ][ 13 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 16 ][ 13 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 17 ][ 13 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 18 ][ 13 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 19 ][ 13 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 20 ][ 13 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 21 ][ 13 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 22 ][ 13 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 23 ][ 13 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 24 ][ 13 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 25 ][ 13 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 0 ][ 12 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 1 ][ 12 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 2 ][ 12 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 3 ][ 12 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 4 ][ 12 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 5 ][ 12 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 6 ][ 12 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 7 ][ 12 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 8 ][ 12 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 9 ][ 12 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 10 ][ 12 ]; 
		 end
		 {1'd1, 5'd17} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 11 ][ 13 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 12 ][ 13 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 13 ][ 13 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 14 ][ 13 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 15 ][ 13 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 16 ][ 13 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 17 ][ 13 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 18 ][ 13 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 19 ][ 13 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 20 ][ 13 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 21 ][ 13 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 22 ][ 13 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 23 ][ 13 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 24 ][ 13 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 25 ][ 13 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 0 ][ 12 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 1 ][ 12 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 2 ][ 12 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 3 ][ 12 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 4 ][ 12 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 5 ][ 12 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 6 ][ 12 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 7 ][ 12 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 8 ][ 12 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 9 ][ 12 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 10 ][ 12 ]; 
		 end
		 {1'd1, 5'd18} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = fifoOut[ 41 ][ 1 ]; 
			 muxOutWire[ 18 ] = fifoOut[ 42 ][ 1 ]; 
			 muxOutWire[ 19 ] = fifoOut[ 43 ][ 1 ]; 
			 muxOutWire[ 20 ] = fifoOut[ 44 ][ 1 ]; 
			 muxOutWire[ 21 ] = fifoOut[ 45 ][ 1 ]; 
			 muxOutWire[ 22 ] = fifoOut[ 46 ][ 1 ]; 
			 muxOutWire[ 23 ] = fifoOut[ 47 ][ 1 ]; 
			 muxOutWire[ 24 ] = fifoOut[ 48 ][ 1 ]; 
			 muxOutWire[ 25 ] = fifoOut[ 49 ][ 1 ]; 
			 muxOutWire[ 26 ] = fifoOut[ 11 ][ 13 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 12 ][ 13 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 13 ][ 13 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 14 ][ 13 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 15 ][ 13 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 16 ][ 13 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 17 ][ 13 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 18 ][ 13 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 19 ][ 13 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 20 ][ 13 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 21 ][ 13 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 22 ][ 13 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 23 ][ 13 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 24 ][ 13 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 25 ][ 13 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 0 ][ 12 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 1 ][ 12 ]; 
			 muxOutWire[ 43 ] = fifoOut[ 2 ][ 12 ]; 
			 muxOutWire[ 44 ] = fifoOut[ 3 ][ 12 ]; 
			 muxOutWire[ 45 ] = fifoOut[ 4 ][ 12 ]; 
			 muxOutWire[ 46 ] = fifoOut[ 5 ][ 12 ]; 
			 muxOutWire[ 47 ] = fifoOut[ 6 ][ 12 ]; 
			 muxOutWire[ 48 ] = fifoOut[ 7 ][ 12 ]; 
			 muxOutWire[ 49 ] = fifoOut[ 8 ][ 12 ]; 
			 muxOutWire[ 50 ] = fifoOut[ 9 ][ 12 ]; 
			 muxOutWire[ 51 ] = fifoOut[ 10 ][ 12 ]; 
		 end
		 {1'd1, 5'd19} : begin 
			 muxOutWire[ 0 ] = fifoOut[ 50 ][ 2 ]; 
			 muxOutWire[ 1 ] = fifoOut[ 51 ][ 2 ]; 
			 muxOutWire[ 2 ] = fifoOut[ 26 ][ 1 ]; 
			 muxOutWire[ 3 ] = fifoOut[ 27 ][ 1 ]; 
			 muxOutWire[ 4 ] = fifoOut[ 28 ][ 1 ]; 
			 muxOutWire[ 5 ] = fifoOut[ 29 ][ 1 ]; 
			 muxOutWire[ 6 ] = fifoOut[ 30 ][ 1 ]; 
			 muxOutWire[ 7 ] = fifoOut[ 31 ][ 1 ]; 
			 muxOutWire[ 8 ] = fifoOut[ 32 ][ 1 ]; 
			 muxOutWire[ 9 ] = fifoOut[ 33 ][ 1 ]; 
			 muxOutWire[ 10 ] = fifoOut[ 34 ][ 1 ]; 
			 muxOutWire[ 11 ] = fifoOut[ 35 ][ 1 ]; 
			 muxOutWire[ 12 ] = fifoOut[ 36 ][ 1 ]; 
			 muxOutWire[ 13 ] = fifoOut[ 37 ][ 1 ]; 
			 muxOutWire[ 14 ] = fifoOut[ 38 ][ 1 ]; 
			 muxOutWire[ 15 ] = fifoOut[ 39 ][ 1 ]; 
			 muxOutWire[ 16 ] = fifoOut[ 40 ][ 1 ]; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = fifoOut[ 11 ][ 13 ]; 
			 muxOutWire[ 27 ] = fifoOut[ 12 ][ 13 ]; 
			 muxOutWire[ 28 ] = fifoOut[ 13 ][ 13 ]; 
			 muxOutWire[ 29 ] = fifoOut[ 14 ][ 13 ]; 
			 muxOutWire[ 30 ] = fifoOut[ 15 ][ 13 ]; 
			 muxOutWire[ 31 ] = fifoOut[ 16 ][ 13 ]; 
			 muxOutWire[ 32 ] = fifoOut[ 17 ][ 13 ]; 
			 muxOutWire[ 33 ] = fifoOut[ 18 ][ 13 ]; 
			 muxOutWire[ 34 ] = fifoOut[ 19 ][ 13 ]; 
			 muxOutWire[ 35 ] = fifoOut[ 20 ][ 13 ]; 
			 muxOutWire[ 36 ] = fifoOut[ 21 ][ 13 ]; 
			 muxOutWire[ 37 ] = fifoOut[ 22 ][ 13 ]; 
			 muxOutWire[ 38 ] = fifoOut[ 23 ][ 13 ]; 
			 muxOutWire[ 39 ] = fifoOut[ 24 ][ 13 ]; 
			 muxOutWire[ 40 ] = fifoOut[ 25 ][ 13 ]; 
			 muxOutWire[ 41 ] = fifoOut[ 0 ][ 12 ]; 
			 muxOutWire[ 42 ] = fifoOut[ 1 ][ 12 ]; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
		 end
    default:begin 
			 muxOutWire[ 0 ] = 0; 
			 muxOutWire[ 1 ] = 0; 
			 muxOutWire[ 2 ] = 0; 
			 muxOutWire[ 3 ] = 0; 
			 muxOutWire[ 4 ] = 0; 
			 muxOutWire[ 5 ] = 0; 
			 muxOutWire[ 6 ] = 0; 
			 muxOutWire[ 7 ] = 0; 
			 muxOutWire[ 8 ] = 0; 
			 muxOutWire[ 9 ] = 0; 
			 muxOutWire[ 10 ] = 0; 
			 muxOutWire[ 11 ] = 0; 
			 muxOutWire[ 12 ] = 0; 
			 muxOutWire[ 13 ] = 0; 
			 muxOutWire[ 14 ] = 0; 
			 muxOutWire[ 15 ] = 0; 
			 muxOutWire[ 16 ] = 0; 
			 muxOutWire[ 17 ] = 0; 
			 muxOutWire[ 18 ] = 0; 
			 muxOutWire[ 19 ] = 0; 
			 muxOutWire[ 20 ] = 0; 
			 muxOutWire[ 21 ] = 0; 
			 muxOutWire[ 22 ] = 0; 
			 muxOutWire[ 23 ] = 0; 
			 muxOutWire[ 24 ] = 0; 
			 muxOutWire[ 25 ] = 0; 
			 muxOutWire[ 26 ] = 0; 
			 muxOutWire[ 27 ] = 0; 
			 muxOutWire[ 28 ] = 0; 
			 muxOutWire[ 29 ] = 0; 
			 muxOutWire[ 30 ] = 0; 
			 muxOutWire[ 31 ] = 0; 
			 muxOutWire[ 32 ] = 0; 
			 muxOutWire[ 33 ] = 0; 
			 muxOutWire[ 34 ] = 0; 
			 muxOutWire[ 35 ] = 0; 
			 muxOutWire[ 36 ] = 0; 
			 muxOutWire[ 37 ] = 0; 
			 muxOutWire[ 38 ] = 0; 
			 muxOutWire[ 39 ] = 0; 
			 muxOutWire[ 40 ] = 0; 
			 muxOutWire[ 41 ] = 0; 
			 muxOutWire[ 42 ] = 0; 
			 muxOutWire[ 43 ] = 0; 
			 muxOutWire[ 44 ] = 0; 
			 muxOutWire[ 45 ] = 0; 
			 muxOutWire[ 46 ] = 0; 
			 muxOutWire[ 47 ] = 0; 
			 muxOutWire[ 48 ] = 0; 
			 muxOutWire[ 49 ] = 0; 
			 muxOutWire[ 50 ] = 0; 
			 muxOutWire[ 51 ] = 0; 
    end
    endcase
end
endmodule
