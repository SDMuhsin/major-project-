`timescale 1ns / 1ps
module LMem1To0_511_circ14_yesshift_nounload_scripted(
        muxOut,
        ly0In,
        wr_en,
        feedback_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 14;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

input feedback_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        if(feedback_en) begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= fifoOut[i][c-1];
         end
        end
        else begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= ly0InConnector[i];
         end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[18][2];
              muxOutConnector[1] = fifoOut[19][2];
              muxOutConnector[2] = fifoOut[20][2];
              muxOutConnector[3] = fifoOut[21][2];
              muxOutConnector[4] = fifoOut[22][2];
              muxOutConnector[5] = fifoOut[23][2];
              muxOutConnector[6] = fifoOut[24][2];
              muxOutConnector[7] = fifoOut[25][2];
              muxOutConnector[8] = fifoOut[0][1];
              muxOutConnector[9] = fifoOut[1][1];
              muxOutConnector[10] = fifoOut[2][1];
              muxOutConnector[11] = fifoOut[3][1];
              muxOutConnector[12] = fifoOut[4][1];
              muxOutConnector[13] = fifoOut[5][1];
              muxOutConnector[14] = fifoOut[6][1];
              muxOutConnector[15] = fifoOut[7][1];
              muxOutConnector[16] = fifoOut[8][1];
              muxOutConnector[17] = fifoOut[9][1];
              muxOutConnector[18] = fifoOut[10][1];
              muxOutConnector[19] = fifoOut[11][1];
              muxOutConnector[20] = fifoOut[12][1];
              muxOutConnector[21] = fifoOut[13][1];
              muxOutConnector[22] = fifoOut[14][1];
              muxOutConnector[23] = fifoOut[15][1];
              muxOutConnector[24] = fifoOut[16][1];
              muxOutConnector[25] = fifoOut[17][1];
              muxOutConnector[26] = fifoOut[14][12];
              muxOutConnector[27] = fifoOut[15][12];
              muxOutConnector[28] = fifoOut[16][12];
              muxOutConnector[29] = fifoOut[17][12];
              muxOutConnector[30] = fifoOut[18][12];
              muxOutConnector[31] = fifoOut[19][12];
              muxOutConnector[32] = fifoOut[20][12];
              muxOutConnector[33] = fifoOut[21][12];
              muxOutConnector[34] = fifoOut[22][12];
              muxOutConnector[35] = fifoOut[23][12];
              muxOutConnector[36] = fifoOut[24][12];
              muxOutConnector[37] = fifoOut[25][12];
              muxOutConnector[38] = fifoOut[0][11];
              muxOutConnector[39] = fifoOut[1][11];
              muxOutConnector[40] = fifoOut[2][11];
              muxOutConnector[41] = fifoOut[3][11];
              muxOutConnector[42] = fifoOut[4][11];
              muxOutConnector[43] = fifoOut[5][11];
              muxOutConnector[44] = fifoOut[6][11];
              muxOutConnector[45] = fifoOut[7][11];
              muxOutConnector[46] = fifoOut[8][11];
              muxOutConnector[47] = fifoOut[9][11];
              muxOutConnector[48] = fifoOut[10][11];
              muxOutConnector[49] = fifoOut[11][11];
              muxOutConnector[50] = fifoOut[12][11];
              muxOutConnector[51] = fifoOut[13][11];
       end
       1: begin
              muxOutConnector[0] = fifoOut[18][2];
              muxOutConnector[1] = fifoOut[19][2];
              muxOutConnector[2] = fifoOut[20][2];
              muxOutConnector[3] = fifoOut[21][2];
              muxOutConnector[4] = fifoOut[22][2];
              muxOutConnector[5] = fifoOut[23][2];
              muxOutConnector[6] = fifoOut[24][2];
              muxOutConnector[7] = fifoOut[25][2];
              muxOutConnector[8] = fifoOut[0][1];
              muxOutConnector[9] = fifoOut[1][1];
              muxOutConnector[10] = fifoOut[2][1];
              muxOutConnector[11] = fifoOut[3][1];
              muxOutConnector[12] = fifoOut[4][1];
              muxOutConnector[13] = fifoOut[5][1];
              muxOutConnector[14] = fifoOut[6][1];
              muxOutConnector[15] = fifoOut[7][1];
              muxOutConnector[16] = fifoOut[8][1];
              muxOutConnector[17] = fifoOut[9][1];
              muxOutConnector[18] = fifoOut[10][1];
              muxOutConnector[19] = fifoOut[11][1];
              muxOutConnector[20] = fifoOut[12][1];
              muxOutConnector[21] = fifoOut[13][1];
              muxOutConnector[22] = fifoOut[14][1];
              muxOutConnector[23] = fifoOut[15][1];
              muxOutConnector[24] = fifoOut[16][1];
              muxOutConnector[25] = fifoOut[50][0];
              muxOutConnector[26] = fifoOut[14][12];
              muxOutConnector[27] = fifoOut[15][12];
              muxOutConnector[28] = fifoOut[16][12];
              muxOutConnector[29] = fifoOut[17][12];
              muxOutConnector[30] = fifoOut[18][12];
              muxOutConnector[31] = fifoOut[19][12];
              muxOutConnector[32] = fifoOut[20][12];
              muxOutConnector[33] = fifoOut[21][12];
              muxOutConnector[34] = fifoOut[22][12];
              muxOutConnector[35] = fifoOut[23][12];
              muxOutConnector[36] = fifoOut[24][12];
              muxOutConnector[37] = fifoOut[25][12];
              muxOutConnector[38] = fifoOut[0][11];
              muxOutConnector[39] = fifoOut[1][11];
              muxOutConnector[40] = fifoOut[2][11];
              muxOutConnector[41] = fifoOut[3][11];
              muxOutConnector[42] = fifoOut[4][11];
              muxOutConnector[43] = fifoOut[5][11];
              muxOutConnector[44] = fifoOut[6][11];
              muxOutConnector[45] = fifoOut[7][11];
              muxOutConnector[46] = fifoOut[8][11];
              muxOutConnector[47] = fifoOut[9][11];
              muxOutConnector[48] = fifoOut[10][11];
              muxOutConnector[49] = fifoOut[11][11];
              muxOutConnector[50] = fifoOut[12][11];
              muxOutConnector[51] = fifoOut[13][11];
       end
       2: begin
              muxOutConnector[0] = fifoOut[51][1];
              muxOutConnector[1] = fifoOut[26][0];
              muxOutConnector[2] = fifoOut[27][0];
              muxOutConnector[3] = fifoOut[28][0];
              muxOutConnector[4] = fifoOut[29][0];
              muxOutConnector[5] = fifoOut[30][0];
              muxOutConnector[6] = fifoOut[31][0];
              muxOutConnector[7] = fifoOut[32][0];
              muxOutConnector[8] = fifoOut[33][0];
              muxOutConnector[9] = fifoOut[34][0];
              muxOutConnector[10] = fifoOut[35][0];
              muxOutConnector[11] = fifoOut[36][0];
              muxOutConnector[12] = fifoOut[37][0];
              muxOutConnector[13] = fifoOut[38][0];
              muxOutConnector[14] = fifoOut[39][0];
              muxOutConnector[15] = fifoOut[40][0];
              muxOutConnector[16] = fifoOut[41][0];
              muxOutConnector[17] = fifoOut[42][0];
              muxOutConnector[18] = fifoOut[43][0];
              muxOutConnector[19] = fifoOut[44][0];
              muxOutConnector[20] = fifoOut[45][0];
              muxOutConnector[21] = fifoOut[46][0];
              muxOutConnector[22] = fifoOut[47][0];
              muxOutConnector[23] = fifoOut[48][0];
              muxOutConnector[24] = fifoOut[49][0];
              muxOutConnector[25] = fifoOut[50][0];
              muxOutConnector[26] = fifoOut[14][12];
              muxOutConnector[27] = fifoOut[15][12];
              muxOutConnector[28] = fifoOut[16][12];
              muxOutConnector[29] = fifoOut[17][12];
              muxOutConnector[30] = fifoOut[18][12];
              muxOutConnector[31] = fifoOut[19][12];
              muxOutConnector[32] = fifoOut[20][12];
              muxOutConnector[33] = fifoOut[21][12];
              muxOutConnector[34] = fifoOut[22][12];
              muxOutConnector[35] = fifoOut[23][12];
              muxOutConnector[36] = fifoOut[24][12];
              muxOutConnector[37] = fifoOut[25][12];
              muxOutConnector[38] = fifoOut[0][11];
              muxOutConnector[39] = fifoOut[1][11];
              muxOutConnector[40] = fifoOut[2][11];
              muxOutConnector[41] = fifoOut[3][11];
              muxOutConnector[42] = fifoOut[4][11];
              muxOutConnector[43] = fifoOut[5][11];
              muxOutConnector[44] = fifoOut[6][11];
              muxOutConnector[45] = fifoOut[7][11];
              muxOutConnector[46] = fifoOut[8][11];
              muxOutConnector[47] = fifoOut[9][11];
              muxOutConnector[48] = fifoOut[10][11];
              muxOutConnector[49] = fifoOut[11][11];
              muxOutConnector[50] = fifoOut[12][11];
              muxOutConnector[51] = fifoOut[13][11];
       end
       3: begin
              muxOutConnector[0] = fifoOut[51][1];
              muxOutConnector[1] = fifoOut[26][0];
              muxOutConnector[2] = fifoOut[27][0];
              muxOutConnector[3] = fifoOut[28][0];
              muxOutConnector[4] = fifoOut[29][0];
              muxOutConnector[5] = fifoOut[30][0];
              muxOutConnector[6] = fifoOut[31][0];
              muxOutConnector[7] = fifoOut[32][0];
              muxOutConnector[8] = fifoOut[33][0];
              muxOutConnector[9] = fifoOut[34][0];
              muxOutConnector[10] = fifoOut[35][0];
              muxOutConnector[11] = fifoOut[36][0];
              muxOutConnector[12] = fifoOut[37][0];
              muxOutConnector[13] = fifoOut[38][0];
              muxOutConnector[14] = fifoOut[39][0];
              muxOutConnector[15] = fifoOut[40][0];
              muxOutConnector[16] = fifoOut[41][0];
              muxOutConnector[17] = fifoOut[42][0];
              muxOutConnector[18] = fifoOut[43][0];
              muxOutConnector[19] = fifoOut[44][0];
              muxOutConnector[20] = fifoOut[45][0];
              muxOutConnector[21] = fifoOut[46][0];
              muxOutConnector[22] = fifoOut[47][0];
              muxOutConnector[23] = fifoOut[48][0];
              muxOutConnector[24] = fifoOut[49][0];
              muxOutConnector[25] = fifoOut[50][0];
              muxOutConnector[26] = fifoOut[14][12];
              muxOutConnector[27] = fifoOut[15][12];
              muxOutConnector[28] = fifoOut[16][12];
              muxOutConnector[29] = fifoOut[17][12];
              muxOutConnector[30] = fifoOut[18][12];
              muxOutConnector[31] = fifoOut[19][12];
              muxOutConnector[32] = fifoOut[20][12];
              muxOutConnector[33] = fifoOut[21][12];
              muxOutConnector[34] = fifoOut[22][12];
              muxOutConnector[35] = fifoOut[23][12];
              muxOutConnector[36] = fifoOut[24][12];
              muxOutConnector[37] = fifoOut[25][12];
              muxOutConnector[38] = fifoOut[0][11];
              muxOutConnector[39] = fifoOut[1][11];
              muxOutConnector[40] = fifoOut[2][11];
              muxOutConnector[41] = fifoOut[3][11];
              muxOutConnector[42] = fifoOut[4][11];
              muxOutConnector[43] = fifoOut[5][11];
              muxOutConnector[44] = fifoOut[6][11];
              muxOutConnector[45] = fifoOut[7][11];
              muxOutConnector[46] = fifoOut[8][11];
              muxOutConnector[47] = fifoOut[9][11];
              muxOutConnector[48] = fifoOut[10][11];
              muxOutConnector[49] = fifoOut[11][11];
              muxOutConnector[50] = fifoOut[12][11];
              muxOutConnector[51] = fifoOut[13][11];
       end
       4: begin
              muxOutConnector[0] = fifoOut[51][1];
              muxOutConnector[1] = fifoOut[26][0];
              muxOutConnector[2] = fifoOut[27][0];
              muxOutConnector[3] = fifoOut[28][0];
              muxOutConnector[4] = fifoOut[29][0];
              muxOutConnector[5] = fifoOut[30][0];
              muxOutConnector[6] = fifoOut[31][0];
              muxOutConnector[7] = fifoOut[32][0];
              muxOutConnector[8] = fifoOut[33][0];
              muxOutConnector[9] = fifoOut[34][0];
              muxOutConnector[10] = fifoOut[35][0];
              muxOutConnector[11] = fifoOut[36][0];
              muxOutConnector[12] = fifoOut[37][0];
              muxOutConnector[13] = fifoOut[38][0];
              muxOutConnector[14] = fifoOut[39][0];
              muxOutConnector[15] = fifoOut[40][0];
              muxOutConnector[16] = fifoOut[41][0];
              muxOutConnector[17] = fifoOut[42][0];
              muxOutConnector[18] = fifoOut[43][0];
              muxOutConnector[19] = fifoOut[44][0];
              muxOutConnector[20] = fifoOut[45][0];
              muxOutConnector[21] = fifoOut[46][0];
              muxOutConnector[22] = fifoOut[47][0];
              muxOutConnector[23] = fifoOut[48][0];
              muxOutConnector[24] = fifoOut[49][0];
              muxOutConnector[25] = fifoOut[50][0];
              muxOutConnector[26] = fifoOut[14][12];
              muxOutConnector[27] = fifoOut[15][12];
              muxOutConnector[28] = fifoOut[16][12];
              muxOutConnector[29] = fifoOut[17][12];
              muxOutConnector[30] = fifoOut[18][12];
              muxOutConnector[31] = fifoOut[19][12];
              muxOutConnector[32] = fifoOut[20][12];
              muxOutConnector[33] = fifoOut[21][12];
              muxOutConnector[34] = fifoOut[22][12];
              muxOutConnector[35] = fifoOut[23][12];
              muxOutConnector[36] = fifoOut[24][12];
              muxOutConnector[37] = fifoOut[25][12];
              muxOutConnector[38] = fifoOut[0][11];
              muxOutConnector[39] = fifoOut[1][11];
              muxOutConnector[40] = fifoOut[2][11];
              muxOutConnector[41] = fifoOut[3][11];
              muxOutConnector[42] = fifoOut[4][11];
              muxOutConnector[43] = fifoOut[5][11];
              muxOutConnector[44] = fifoOut[6][11];
              muxOutConnector[45] = fifoOut[7][11];
              muxOutConnector[46] = fifoOut[8][11];
              muxOutConnector[47] = fifoOut[9][11];
              muxOutConnector[48] = fifoOut[10][11];
              muxOutConnector[49] = fifoOut[11][11];
              muxOutConnector[50] = fifoOut[12][11];
              muxOutConnector[51] = fifoOut[13][11];
       end
       5: begin
              muxOutConnector[0] = fifoOut[51][1];
              muxOutConnector[1] = fifoOut[26][0];
              muxOutConnector[2] = fifoOut[27][0];
              muxOutConnector[3] = fifoOut[28][0];
              muxOutConnector[4] = fifoOut[29][0];
              muxOutConnector[5] = fifoOut[30][0];
              muxOutConnector[6] = fifoOut[31][0];
              muxOutConnector[7] = fifoOut[32][0];
              muxOutConnector[8] = fifoOut[33][0];
              muxOutConnector[9] = fifoOut[34][0];
              muxOutConnector[10] = fifoOut[35][0];
              muxOutConnector[11] = fifoOut[36][0];
              muxOutConnector[12] = fifoOut[37][0];
              muxOutConnector[13] = fifoOut[38][0];
              muxOutConnector[14] = fifoOut[39][0];
              muxOutConnector[15] = fifoOut[40][0];
              muxOutConnector[16] = fifoOut[41][0];
              muxOutConnector[17] = fifoOut[42][0];
              muxOutConnector[18] = fifoOut[43][0];
              muxOutConnector[19] = fifoOut[44][0];
              muxOutConnector[20] = fifoOut[45][0];
              muxOutConnector[21] = fifoOut[46][0];
              muxOutConnector[22] = fifoOut[47][0];
              muxOutConnector[23] = fifoOut[48][0];
              muxOutConnector[24] = fifoOut[49][0];
              muxOutConnector[25] = fifoOut[50][0];
              muxOutConnector[26] = fifoOut[14][12];
              muxOutConnector[27] = fifoOut[15][12];
              muxOutConnector[28] = fifoOut[16][12];
              muxOutConnector[29] = fifoOut[17][12];
              muxOutConnector[30] = fifoOut[18][12];
              muxOutConnector[31] = fifoOut[19][12];
              muxOutConnector[32] = fifoOut[20][12];
              muxOutConnector[33] = fifoOut[21][12];
              muxOutConnector[34] = fifoOut[22][12];
              muxOutConnector[35] = fifoOut[23][12];
              muxOutConnector[36] = fifoOut[24][12];
              muxOutConnector[37] = fifoOut[25][12];
              muxOutConnector[38] = fifoOut[0][11];
              muxOutConnector[39] = fifoOut[1][11];
              muxOutConnector[40] = fifoOut[2][11];
              muxOutConnector[41] = fifoOut[3][11];
              muxOutConnector[42] = fifoOut[4][11];
              muxOutConnector[43] = fifoOut[5][11];
              muxOutConnector[44] = fifoOut[6][11];
              muxOutConnector[45] = fifoOut[7][11];
              muxOutConnector[46] = fifoOut[8][11];
              muxOutConnector[47] = fifoOut[9][11];
              muxOutConnector[48] = fifoOut[10][11];
              muxOutConnector[49] = fifoOut[11][11];
              muxOutConnector[50] = fifoOut[12][11];
              muxOutConnector[51] = fifoOut[13][11];
       end
       6: begin
              muxOutConnector[0] = fifoOut[51][1];
              muxOutConnector[1] = fifoOut[26][0];
              muxOutConnector[2] = fifoOut[27][0];
              muxOutConnector[3] = fifoOut[28][0];
              muxOutConnector[4] = fifoOut[29][0];
              muxOutConnector[5] = fifoOut[30][0];
              muxOutConnector[6] = fifoOut[31][0];
              muxOutConnector[7] = fifoOut[32][0];
              muxOutConnector[8] = fifoOut[33][0];
              muxOutConnector[9] = fifoOut[34][0];
              muxOutConnector[10] = fifoOut[35][0];
              muxOutConnector[11] = fifoOut[36][0];
              muxOutConnector[12] = fifoOut[37][0];
              muxOutConnector[13] = fifoOut[38][0];
              muxOutConnector[14] = fifoOut[39][0];
              muxOutConnector[15] = fifoOut[40][0];
              muxOutConnector[16] = fifoOut[41][0];
              muxOutConnector[17] = fifoOut[42][0];
              muxOutConnector[18] = fifoOut[43][0];
              muxOutConnector[19] = fifoOut[44][0];
              muxOutConnector[20] = fifoOut[45][0];
              muxOutConnector[21] = fifoOut[46][0];
              muxOutConnector[22] = fifoOut[47][0];
              muxOutConnector[23] = fifoOut[48][0];
              muxOutConnector[24] = fifoOut[49][0];
              muxOutConnector[25] = fifoOut[50][0];
              muxOutConnector[26] = fifoOut[14][12];
              muxOutConnector[27] = fifoOut[15][12];
              muxOutConnector[28] = fifoOut[16][12];
              muxOutConnector[29] = fifoOut[17][12];
              muxOutConnector[30] = fifoOut[18][12];
              muxOutConnector[31] = fifoOut[19][12];
              muxOutConnector[32] = fifoOut[20][12];
              muxOutConnector[33] = fifoOut[21][12];
              muxOutConnector[34] = fifoOut[22][12];
              muxOutConnector[35] = fifoOut[23][12];
              muxOutConnector[36] = fifoOut[24][12];
              muxOutConnector[37] = fifoOut[25][12];
              muxOutConnector[38] = fifoOut[0][11];
              muxOutConnector[39] = fifoOut[1][11];
              muxOutConnector[40] = fifoOut[2][11];
              muxOutConnector[41] = fifoOut[3][11];
              muxOutConnector[42] = fifoOut[4][11];
              muxOutConnector[43] = fifoOut[5][11];
              muxOutConnector[44] = fifoOut[6][11];
              muxOutConnector[45] = fifoOut[7][11];
              muxOutConnector[46] = fifoOut[8][11];
              muxOutConnector[47] = fifoOut[9][11];
              muxOutConnector[48] = fifoOut[10][11];
              muxOutConnector[49] = fifoOut[11][11];
              muxOutConnector[50] = fifoOut[12][11];
              muxOutConnector[51] = fifoOut[13][11];
       end
       7: begin
              muxOutConnector[0] = fifoOut[51][1];
              muxOutConnector[1] = fifoOut[26][0];
              muxOutConnector[2] = fifoOut[27][0];
              muxOutConnector[3] = fifoOut[28][0];
              muxOutConnector[4] = fifoOut[29][0];
              muxOutConnector[5] = fifoOut[30][0];
              muxOutConnector[6] = fifoOut[31][0];
              muxOutConnector[7] = fifoOut[32][0];
              muxOutConnector[8] = fifoOut[33][0];
              muxOutConnector[9] = fifoOut[34][0];
              muxOutConnector[10] = fifoOut[35][0];
              muxOutConnector[11] = fifoOut[36][0];
              muxOutConnector[12] = fifoOut[37][0];
              muxOutConnector[13] = fifoOut[38][0];
              muxOutConnector[14] = fifoOut[39][0];
              muxOutConnector[15] = fifoOut[40][0];
              muxOutConnector[16] = fifoOut[41][0];
              muxOutConnector[17] = fifoOut[42][0];
              muxOutConnector[18] = fifoOut[43][0];
              muxOutConnector[19] = fifoOut[44][0];
              muxOutConnector[20] = fifoOut[45][0];
              muxOutConnector[21] = fifoOut[46][0];
              muxOutConnector[22] = fifoOut[47][0];
              muxOutConnector[23] = fifoOut[48][0];
              muxOutConnector[24] = fifoOut[49][0];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[14][12];
              muxOutConnector[27] = fifoOut[15][12];
              muxOutConnector[28] = fifoOut[16][12];
              muxOutConnector[29] = fifoOut[17][12];
              muxOutConnector[30] = fifoOut[18][12];
              muxOutConnector[31] = fifoOut[19][12];
              muxOutConnector[32] = fifoOut[20][12];
              muxOutConnector[33] = fifoOut[21][12];
              muxOutConnector[34] = fifoOut[22][12];
              muxOutConnector[35] = fifoOut[23][12];
              muxOutConnector[36] = fifoOut[24][12];
              muxOutConnector[37] = fifoOut[25][12];
              muxOutConnector[38] = fifoOut[0][11];
              muxOutConnector[39] = fifoOut[1][11];
              muxOutConnector[40] = fifoOut[2][11];
              muxOutConnector[41] = fifoOut[3][11];
              muxOutConnector[42] = fifoOut[4][11];
              muxOutConnector[43] = fifoOut[5][11];
              muxOutConnector[44] = fifoOut[6][11];
              muxOutConnector[45] = fifoOut[7][11];
              muxOutConnector[46] = fifoOut[8][11];
              muxOutConnector[47] = fifoOut[9][11];
              muxOutConnector[48] = fifoOut[10][11];
              muxOutConnector[49] = fifoOut[11][11];
              muxOutConnector[50] = fifoOut[12][11];
              muxOutConnector[51] = fifoOut[13][11];
       end
       8: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[14][12];
              muxOutConnector[27] = fifoOut[15][12];
              muxOutConnector[28] = fifoOut[16][12];
              muxOutConnector[29] = fifoOut[17][12];
              muxOutConnector[30] = fifoOut[18][12];
              muxOutConnector[31] = fifoOut[19][12];
              muxOutConnector[32] = fifoOut[20][12];
              muxOutConnector[33] = fifoOut[21][12];
              muxOutConnector[34] = fifoOut[22][12];
              muxOutConnector[35] = fifoOut[23][12];
              muxOutConnector[36] = fifoOut[24][12];
              muxOutConnector[37] = fifoOut[25][12];
              muxOutConnector[38] = fifoOut[0][11];
              muxOutConnector[39] = fifoOut[1][11];
              muxOutConnector[40] = fifoOut[2][11];
              muxOutConnector[41] = fifoOut[3][11];
              muxOutConnector[42] = fifoOut[4][11];
              muxOutConnector[43] = fifoOut[5][11];
              muxOutConnector[44] = fifoOut[6][11];
              muxOutConnector[45] = fifoOut[7][11];
              muxOutConnector[46] = fifoOut[8][11];
              muxOutConnector[47] = fifoOut[9][11];
              muxOutConnector[48] = fifoOut[10][11];
              muxOutConnector[49] = fifoOut[11][11];
              muxOutConnector[50] = fifoOut[12][11];
              muxOutConnector[51] = fifoOut[13][11];
       end
       9: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[14][12];
              muxOutConnector[27] = fifoOut[15][12];
              muxOutConnector[28] = fifoOut[16][12];
              muxOutConnector[29] = fifoOut[17][12];
              muxOutConnector[30] = fifoOut[18][12];
              muxOutConnector[31] = fifoOut[19][12];
              muxOutConnector[32] = fifoOut[20][12];
              muxOutConnector[33] = fifoOut[21][12];
              muxOutConnector[34] = fifoOut[22][12];
              muxOutConnector[35] = fifoOut[23][12];
              muxOutConnector[36] = fifoOut[24][12];
              muxOutConnector[37] = fifoOut[25][12];
              muxOutConnector[38] = fifoOut[0][11];
              muxOutConnector[39] = fifoOut[1][11];
              muxOutConnector[40] = fifoOut[2][11];
              muxOutConnector[41] = fifoOut[3][11];
              muxOutConnector[42] = fifoOut[4][11];
              muxOutConnector[43] = fifoOut[5][11];
              muxOutConnector[44] = fifoOut[6][11];
              muxOutConnector[45] = fifoOut[7][11];
              muxOutConnector[46] = fifoOut[8][11];
              muxOutConnector[47] = fifoOut[9][11];
              muxOutConnector[48] = fifoOut[10][11];
              muxOutConnector[49] = fifoOut[11][11];
              muxOutConnector[50] = fifoOut[12][11];
              muxOutConnector[51] = fifoOut[13][11];
       end
       10: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[14][12];
              muxOutConnector[27] = fifoOut[15][12];
              muxOutConnector[28] = fifoOut[16][12];
              muxOutConnector[29] = fifoOut[17][12];
              muxOutConnector[30] = fifoOut[18][12];
              muxOutConnector[31] = fifoOut[19][12];
              muxOutConnector[32] = fifoOut[20][12];
              muxOutConnector[33] = fifoOut[21][12];
              muxOutConnector[34] = fifoOut[22][12];
              muxOutConnector[35] = fifoOut[23][12];
              muxOutConnector[36] = fifoOut[24][12];
              muxOutConnector[37] = fifoOut[25][12];
              muxOutConnector[38] = fifoOut[0][11];
              muxOutConnector[39] = fifoOut[1][11];
              muxOutConnector[40] = fifoOut[2][11];
              muxOutConnector[41] = fifoOut[3][11];
              muxOutConnector[42] = fifoOut[4][11];
              muxOutConnector[43] = fifoOut[5][11];
              muxOutConnector[44] = fifoOut[6][11];
              muxOutConnector[45] = fifoOut[7][11];
              muxOutConnector[46] = fifoOut[8][11];
              muxOutConnector[47] = fifoOut[9][11];
              muxOutConnector[48] = fifoOut[10][11];
              muxOutConnector[49] = fifoOut[11][11];
              muxOutConnector[50] = fifoOut[12][11];
              muxOutConnector[51] = fifoOut[13][11];
       end
       11: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[14][12];
              muxOutConnector[27] = fifoOut[15][12];
              muxOutConnector[28] = fifoOut[16][12];
              muxOutConnector[29] = fifoOut[17][12];
              muxOutConnector[30] = fifoOut[18][12];
              muxOutConnector[31] = fifoOut[19][12];
              muxOutConnector[32] = fifoOut[20][12];
              muxOutConnector[33] = fifoOut[21][12];
              muxOutConnector[34] = fifoOut[22][12];
              muxOutConnector[35] = fifoOut[23][12];
              muxOutConnector[36] = fifoOut[24][12];
              muxOutConnector[37] = fifoOut[25][12];
              muxOutConnector[38] = fifoOut[0][11];
              muxOutConnector[39] = fifoOut[1][11];
              muxOutConnector[40] = fifoOut[2][11];
              muxOutConnector[41] = fifoOut[3][11];
              muxOutConnector[42] = fifoOut[4][11];
              muxOutConnector[43] = fifoOut[5][11];
              muxOutConnector[44] = fifoOut[6][11];
              muxOutConnector[45] = fifoOut[7][11];
              muxOutConnector[46] = fifoOut[8][11];
              muxOutConnector[47] = fifoOut[9][11];
              muxOutConnector[48] = fifoOut[10][11];
              muxOutConnector[49] = fifoOut[11][11];
              muxOutConnector[50] = fifoOut[12][11];
              muxOutConnector[51] = fifoOut[13][11];
       end
       12: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[14][12];
              muxOutConnector[27] = fifoOut[15][12];
              muxOutConnector[28] = fifoOut[16][12];
              muxOutConnector[29] = fifoOut[50][11];
              muxOutConnector[30] = fifoOut[51][11];
              muxOutConnector[31] = fifoOut[26][10];
              muxOutConnector[32] = fifoOut[27][10];
              muxOutConnector[33] = fifoOut[28][10];
              muxOutConnector[34] = fifoOut[29][10];
              muxOutConnector[35] = fifoOut[30][10];
              muxOutConnector[36] = fifoOut[31][10];
              muxOutConnector[37] = fifoOut[32][10];
              muxOutConnector[38] = fifoOut[33][10];
              muxOutConnector[39] = fifoOut[34][10];
              muxOutConnector[40] = fifoOut[35][10];
              muxOutConnector[41] = fifoOut[36][10];
              muxOutConnector[42] = fifoOut[37][10];
              muxOutConnector[43] = fifoOut[38][10];
              muxOutConnector[44] = fifoOut[39][10];
              muxOutConnector[45] = fifoOut[40][10];
              muxOutConnector[46] = fifoOut[41][10];
              muxOutConnector[47] = fifoOut[42][10];
              muxOutConnector[48] = fifoOut[43][10];
              muxOutConnector[49] = fifoOut[44][10];
              muxOutConnector[50] = fifoOut[45][10];
              muxOutConnector[51] = fifoOut[46][10];
       end
       13: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[47][11];
              muxOutConnector[27] = fifoOut[48][11];
              muxOutConnector[28] = fifoOut[49][11];
              muxOutConnector[29] = fifoOut[50][11];
              muxOutConnector[30] = fifoOut[51][11];
              muxOutConnector[31] = fifoOut[26][10];
              muxOutConnector[32] = fifoOut[27][10];
              muxOutConnector[33] = fifoOut[28][10];
              muxOutConnector[34] = fifoOut[29][10];
              muxOutConnector[35] = fifoOut[30][10];
              muxOutConnector[36] = fifoOut[31][10];
              muxOutConnector[37] = fifoOut[32][10];
              muxOutConnector[38] = fifoOut[33][10];
              muxOutConnector[39] = fifoOut[34][10];
              muxOutConnector[40] = fifoOut[35][10];
              muxOutConnector[41] = fifoOut[36][10];
              muxOutConnector[42] = fifoOut[37][10];
              muxOutConnector[43] = fifoOut[38][10];
              muxOutConnector[44] = fifoOut[39][10];
              muxOutConnector[45] = fifoOut[40][10];
              muxOutConnector[46] = fifoOut[41][10];
              muxOutConnector[47] = fifoOut[42][10];
              muxOutConnector[48] = fifoOut[43][10];
              muxOutConnector[49] = fifoOut[44][10];
              muxOutConnector[50] = fifoOut[45][10];
              muxOutConnector[51] = fifoOut[46][10];
       end
       14: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[47][11];
              muxOutConnector[27] = fifoOut[48][11];
              muxOutConnector[28] = fifoOut[49][11];
              muxOutConnector[29] = fifoOut[50][11];
              muxOutConnector[30] = fifoOut[51][11];
              muxOutConnector[31] = fifoOut[26][10];
              muxOutConnector[32] = fifoOut[27][10];
              muxOutConnector[33] = fifoOut[28][10];
              muxOutConnector[34] = fifoOut[29][10];
              muxOutConnector[35] = fifoOut[30][10];
              muxOutConnector[36] = fifoOut[31][10];
              muxOutConnector[37] = fifoOut[32][10];
              muxOutConnector[38] = fifoOut[33][10];
              muxOutConnector[39] = fifoOut[34][10];
              muxOutConnector[40] = fifoOut[35][10];
              muxOutConnector[41] = fifoOut[36][10];
              muxOutConnector[42] = fifoOut[37][10];
              muxOutConnector[43] = fifoOut[38][10];
              muxOutConnector[44] = fifoOut[39][10];
              muxOutConnector[45] = fifoOut[40][10];
              muxOutConnector[46] = fifoOut[41][10];
              muxOutConnector[47] = fifoOut[42][10];
              muxOutConnector[48] = fifoOut[43][10];
              muxOutConnector[49] = fifoOut[44][10];
              muxOutConnector[50] = fifoOut[45][10];
              muxOutConnector[51] = fifoOut[46][10];
       end
       15: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[47][11];
              muxOutConnector[27] = fifoOut[48][11];
              muxOutConnector[28] = fifoOut[49][11];
              muxOutConnector[29] = fifoOut[50][11];
              muxOutConnector[30] = fifoOut[51][11];
              muxOutConnector[31] = fifoOut[26][10];
              muxOutConnector[32] = fifoOut[27][10];
              muxOutConnector[33] = fifoOut[28][10];
              muxOutConnector[34] = fifoOut[29][10];
              muxOutConnector[35] = fifoOut[30][10];
              muxOutConnector[36] = fifoOut[31][10];
              muxOutConnector[37] = fifoOut[32][10];
              muxOutConnector[38] = fifoOut[33][10];
              muxOutConnector[39] = fifoOut[34][10];
              muxOutConnector[40] = fifoOut[35][10];
              muxOutConnector[41] = fifoOut[36][10];
              muxOutConnector[42] = fifoOut[37][10];
              muxOutConnector[43] = fifoOut[38][10];
              muxOutConnector[44] = fifoOut[39][10];
              muxOutConnector[45] = fifoOut[40][10];
              muxOutConnector[46] = fifoOut[41][10];
              muxOutConnector[47] = fifoOut[42][10];
              muxOutConnector[48] = fifoOut[43][10];
              muxOutConnector[49] = fifoOut[44][10];
              muxOutConnector[50] = fifoOut[45][10];
              muxOutConnector[51] = fifoOut[46][10];
       end
       16: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[47][11];
              muxOutConnector[27] = fifoOut[48][11];
              muxOutConnector[28] = fifoOut[49][11];
              muxOutConnector[29] = fifoOut[50][11];
              muxOutConnector[30] = fifoOut[51][11];
              muxOutConnector[31] = fifoOut[26][10];
              muxOutConnector[32] = fifoOut[27][10];
              muxOutConnector[33] = fifoOut[28][10];
              muxOutConnector[34] = fifoOut[29][10];
              muxOutConnector[35] = fifoOut[30][10];
              muxOutConnector[36] = fifoOut[31][10];
              muxOutConnector[37] = fifoOut[32][10];
              muxOutConnector[38] = fifoOut[33][10];
              muxOutConnector[39] = fifoOut[34][10];
              muxOutConnector[40] = fifoOut[35][10];
              muxOutConnector[41] = fifoOut[36][10];
              muxOutConnector[42] = fifoOut[37][10];
              muxOutConnector[43] = fifoOut[38][10];
              muxOutConnector[44] = fifoOut[39][10];
              muxOutConnector[45] = fifoOut[40][10];
              muxOutConnector[46] = fifoOut[41][10];
              muxOutConnector[47] = fifoOut[42][10];
              muxOutConnector[48] = fifoOut[43][10];
              muxOutConnector[49] = fifoOut[44][10];
              muxOutConnector[50] = fifoOut[45][10];
              muxOutConnector[51] = fifoOut[46][10];
       end
       17: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[47][11];
              muxOutConnector[27] = fifoOut[48][11];
              muxOutConnector[28] = fifoOut[49][11];
              muxOutConnector[29] = fifoOut[50][11];
              muxOutConnector[30] = fifoOut[51][11];
              muxOutConnector[31] = fifoOut[26][10];
              muxOutConnector[32] = fifoOut[27][10];
              muxOutConnector[33] = fifoOut[28][10];
              muxOutConnector[34] = fifoOut[29][10];
              muxOutConnector[35] = fifoOut[30][10];
              muxOutConnector[36] = fifoOut[31][10];
              muxOutConnector[37] = fifoOut[32][10];
              muxOutConnector[38] = fifoOut[33][10];
              muxOutConnector[39] = fifoOut[34][10];
              muxOutConnector[40] = fifoOut[35][10];
              muxOutConnector[41] = fifoOut[36][10];
              muxOutConnector[42] = fifoOut[37][10];
              muxOutConnector[43] = fifoOut[38][10];
              muxOutConnector[44] = fifoOut[39][10];
              muxOutConnector[45] = fifoOut[40][10];
              muxOutConnector[46] = fifoOut[41][10];
              muxOutConnector[47] = fifoOut[42][10];
              muxOutConnector[48] = fifoOut[43][10];
              muxOutConnector[49] = fifoOut[44][10];
              muxOutConnector[50] = fifoOut[45][10];
              muxOutConnector[51] = fifoOut[46][10];
       end
       18: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[47][11];
              muxOutConnector[27] = fifoOut[48][11];
              muxOutConnector[28] = fifoOut[49][11];
              muxOutConnector[29] = fifoOut[50][11];
              muxOutConnector[30] = fifoOut[51][11];
              muxOutConnector[31] = fifoOut[26][10];
              muxOutConnector[32] = fifoOut[27][10];
              muxOutConnector[33] = fifoOut[28][10];
              muxOutConnector[34] = fifoOut[29][10];
              muxOutConnector[35] = fifoOut[30][10];
              muxOutConnector[36] = fifoOut[31][10];
              muxOutConnector[37] = fifoOut[32][10];
              muxOutConnector[38] = fifoOut[33][10];
              muxOutConnector[39] = fifoOut[34][10];
              muxOutConnector[40] = fifoOut[35][10];
              muxOutConnector[41] = fifoOut[36][10];
              muxOutConnector[42] = fifoOut[37][10];
              muxOutConnector[43] = fifoOut[38][10];
              muxOutConnector[44] = fifoOut[39][10];
              muxOutConnector[45] = fifoOut[40][10];
              muxOutConnector[46] = fifoOut[41][10];
              muxOutConnector[47] = fifoOut[42][10];
              muxOutConnector[48] = fifoOut[43][10];
              muxOutConnector[49] = fifoOut[44][10];
              muxOutConnector[50] = fifoOut[45][10];
              muxOutConnector[51] = fifoOut[46][10];
       end
       19: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[47][11];
              muxOutConnector[27] = fifoOut[48][11];
              muxOutConnector[28] = fifoOut[49][11];
              muxOutConnector[29] = fifoOut[50][11];
              muxOutConnector[30] = fifoOut[51][11];
              muxOutConnector[31] = fifoOut[26][10];
              muxOutConnector[32] = fifoOut[27][10];
              muxOutConnector[33] = fifoOut[28][10];
              muxOutConnector[34] = fifoOut[29][10];
              muxOutConnector[35] = fifoOut[30][10];
              muxOutConnector[36] = fifoOut[31][10];
              muxOutConnector[37] = fifoOut[32][10];
              muxOutConnector[38] = fifoOut[33][10];
              muxOutConnector[39] = fifoOut[34][10];
              muxOutConnector[40] = fifoOut[35][10];
              muxOutConnector[41] = fifoOut[36][10];
              muxOutConnector[42] = fifoOut[37][10];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
