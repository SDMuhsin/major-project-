`timescale 1ns / 1ps
module LMem1To0_511_circ10_yesshift_nounload_scripted(
        muxOut,
        ly0In,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 12;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            fifoOut[i][0] <= ly0InConnector[i];
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[25][4];
              muxOutConnector[1] = fifoOut[0][3];
              muxOutConnector[2] = fifoOut[1][3];
              muxOutConnector[3] = fifoOut[2][3];
              muxOutConnector[4] = fifoOut[3][3];
              muxOutConnector[5] = fifoOut[4][3];
              muxOutConnector[6] = fifoOut[5][3];
              muxOutConnector[7] = fifoOut[6][3];
              muxOutConnector[8] = fifoOut[7][3];
              muxOutConnector[9] = fifoOut[8][3];
              muxOutConnector[10] = fifoOut[9][3];
              muxOutConnector[11] = fifoOut[10][3];
              muxOutConnector[12] = fifoOut[11][3];
              muxOutConnector[13] = fifoOut[12][3];
              muxOutConnector[14] = fifoOut[13][3];
              muxOutConnector[15] = fifoOut[14][3];
              muxOutConnector[16] = fifoOut[15][3];
              muxOutConnector[17] = fifoOut[16][3];
              muxOutConnector[18] = fifoOut[17][3];
              muxOutConnector[19] = fifoOut[18][3];
              muxOutConnector[20] = fifoOut[19][3];
              muxOutConnector[21] = fifoOut[20][3];
              muxOutConnector[22] = fifoOut[21][3];
              muxOutConnector[23] = fifoOut[22][3];
              muxOutConnector[24] = fifoOut[23][3];
              muxOutConnector[25] = fifoOut[24][3];
              muxOutConnector[26] = fifoOut[27][6];
              muxOutConnector[27] = fifoOut[28][6];
              muxOutConnector[28] = fifoOut[29][6];
              muxOutConnector[29] = fifoOut[30][6];
              muxOutConnector[30] = fifoOut[31][6];
              muxOutConnector[31] = fifoOut[32][6];
              muxOutConnector[32] = fifoOut[33][6];
              muxOutConnector[33] = fifoOut[34][6];
              muxOutConnector[34] = fifoOut[35][6];
              muxOutConnector[35] = fifoOut[36][6];
              muxOutConnector[36] = fifoOut[37][6];
              muxOutConnector[37] = fifoOut[38][6];
              muxOutConnector[38] = fifoOut[39][6];
              muxOutConnector[39] = fifoOut[40][6];
              muxOutConnector[40] = fifoOut[41][6];
              muxOutConnector[41] = fifoOut[42][6];
              muxOutConnector[42] = fifoOut[43][6];
              muxOutConnector[43] = fifoOut[44][6];
              muxOutConnector[44] = fifoOut[45][6];
              muxOutConnector[45] = fifoOut[46][6];
              muxOutConnector[46] = fifoOut[47][6];
              muxOutConnector[47] = fifoOut[48][6];
              muxOutConnector[48] = fifoOut[49][6];
              muxOutConnector[49] = fifoOut[50][6];
              muxOutConnector[50] = fifoOut[51][6];
              muxOutConnector[51] = fifoOut[26][5];
       end
       1: begin
              muxOutConnector[0] = fifoOut[25][4];
              muxOutConnector[1] = fifoOut[0][3];
              muxOutConnector[2] = fifoOut[1][3];
              muxOutConnector[3] = fifoOut[2][3];
              muxOutConnector[4] = fifoOut[3][3];
              muxOutConnector[5] = fifoOut[4][3];
              muxOutConnector[6] = fifoOut[5][3];
              muxOutConnector[7] = fifoOut[6][3];
              muxOutConnector[8] = fifoOut[7][3];
              muxOutConnector[9] = fifoOut[8][3];
              muxOutConnector[10] = fifoOut[9][3];
              muxOutConnector[11] = fifoOut[10][3];
              muxOutConnector[12] = fifoOut[11][3];
              muxOutConnector[13] = fifoOut[12][3];
              muxOutConnector[14] = fifoOut[13][3];
              muxOutConnector[15] = fifoOut[14][3];
              muxOutConnector[16] = fifoOut[15][3];
              muxOutConnector[17] = fifoOut[16][3];
              muxOutConnector[18] = fifoOut[17][3];
              muxOutConnector[19] = fifoOut[18][3];
              muxOutConnector[20] = fifoOut[19][3];
              muxOutConnector[21] = fifoOut[20][3];
              muxOutConnector[22] = fifoOut[21][3];
              muxOutConnector[23] = fifoOut[22][3];
              muxOutConnector[24] = fifoOut[23][3];
              muxOutConnector[25] = fifoOut[24][3];
              muxOutConnector[26] = fifoOut[27][6];
              muxOutConnector[27] = fifoOut[28][6];
              muxOutConnector[28] = fifoOut[29][6];
              muxOutConnector[29] = fifoOut[30][6];
              muxOutConnector[30] = fifoOut[31][6];
              muxOutConnector[31] = fifoOut[32][6];
              muxOutConnector[32] = fifoOut[33][6];
              muxOutConnector[33] = fifoOut[34][6];
              muxOutConnector[34] = fifoOut[35][6];
              muxOutConnector[35] = fifoOut[36][6];
              muxOutConnector[36] = fifoOut[37][6];
              muxOutConnector[37] = fifoOut[38][6];
              muxOutConnector[38] = fifoOut[39][6];
              muxOutConnector[39] = fifoOut[40][6];
              muxOutConnector[40] = fifoOut[41][6];
              muxOutConnector[41] = fifoOut[42][6];
              muxOutConnector[42] = fifoOut[43][6];
              muxOutConnector[43] = fifoOut[44][6];
              muxOutConnector[44] = fifoOut[45][6];
              muxOutConnector[45] = fifoOut[46][6];
              muxOutConnector[46] = fifoOut[47][6];
              muxOutConnector[47] = fifoOut[48][6];
              muxOutConnector[48] = fifoOut[49][6];
              muxOutConnector[49] = fifoOut[50][6];
              muxOutConnector[50] = fifoOut[51][6];
              muxOutConnector[51] = fifoOut[26][5];
       end
       2: begin
              muxOutConnector[0] = fifoOut[25][4];
              muxOutConnector[1] = fifoOut[0][3];
              muxOutConnector[2] = fifoOut[1][3];
              muxOutConnector[3] = fifoOut[2][3];
              muxOutConnector[4] = fifoOut[3][3];
              muxOutConnector[5] = fifoOut[4][3];
              muxOutConnector[6] = fifoOut[5][3];
              muxOutConnector[7] = fifoOut[6][3];
              muxOutConnector[8] = fifoOut[7][3];
              muxOutConnector[9] = fifoOut[8][3];
              muxOutConnector[10] = fifoOut[9][3];
              muxOutConnector[11] = fifoOut[10][3];
              muxOutConnector[12] = fifoOut[11][3];
              muxOutConnector[13] = fifoOut[12][3];
              muxOutConnector[14] = fifoOut[13][3];
              muxOutConnector[15] = fifoOut[14][3];
              muxOutConnector[16] = fifoOut[15][3];
              muxOutConnector[17] = fifoOut[16][3];
              muxOutConnector[18] = fifoOut[17][3];
              muxOutConnector[19] = fifoOut[18][3];
              muxOutConnector[20] = fifoOut[19][3];
              muxOutConnector[21] = fifoOut[20][3];
              muxOutConnector[22] = fifoOut[21][3];
              muxOutConnector[23] = fifoOut[22][3];
              muxOutConnector[24] = fifoOut[23][3];
              muxOutConnector[25] = fifoOut[24][3];
              muxOutConnector[26] = fifoOut[27][6];
              muxOutConnector[27] = fifoOut[28][6];
              muxOutConnector[28] = fifoOut[29][6];
              muxOutConnector[29] = fifoOut[30][6];
              muxOutConnector[30] = fifoOut[31][6];
              muxOutConnector[31] = fifoOut[32][6];
              muxOutConnector[32] = fifoOut[33][6];
              muxOutConnector[33] = fifoOut[34][6];
              muxOutConnector[34] = fifoOut[35][6];
              muxOutConnector[35] = fifoOut[36][6];
              muxOutConnector[36] = fifoOut[37][6];
              muxOutConnector[37] = fifoOut[38][6];
              muxOutConnector[38] = fifoOut[39][6];
              muxOutConnector[39] = fifoOut[40][6];
              muxOutConnector[40] = fifoOut[41][6];
              muxOutConnector[41] = fifoOut[42][6];
              muxOutConnector[42] = fifoOut[43][6];
              muxOutConnector[43] = fifoOut[44][6];
              muxOutConnector[44] = fifoOut[45][6];
              muxOutConnector[45] = fifoOut[46][6];
              muxOutConnector[46] = fifoOut[47][6];
              muxOutConnector[47] = fifoOut[48][6];
              muxOutConnector[48] = fifoOut[49][6];
              muxOutConnector[49] = fifoOut[50][6];
              muxOutConnector[50] = fifoOut[51][6];
              muxOutConnector[51] = fifoOut[26][5];
       end
       3: begin
              muxOutConnector[0] = fifoOut[25][4];
              muxOutConnector[1] = fifoOut[0][3];
              muxOutConnector[2] = fifoOut[1][3];
              muxOutConnector[3] = fifoOut[2][3];
              muxOutConnector[4] = fifoOut[3][3];
              muxOutConnector[5] = fifoOut[4][3];
              muxOutConnector[6] = fifoOut[5][3];
              muxOutConnector[7] = fifoOut[6][3];
              muxOutConnector[8] = fifoOut[7][3];
              muxOutConnector[9] = fifoOut[8][3];
              muxOutConnector[10] = fifoOut[9][3];
              muxOutConnector[11] = fifoOut[10][3];
              muxOutConnector[12] = fifoOut[11][3];
              muxOutConnector[13] = fifoOut[12][3];
              muxOutConnector[14] = fifoOut[13][3];
              muxOutConnector[15] = fifoOut[14][3];
              muxOutConnector[16] = fifoOut[15][3];
              muxOutConnector[17] = fifoOut[16][3];
              muxOutConnector[18] = fifoOut[46][2];
              muxOutConnector[19] = fifoOut[47][2];
              muxOutConnector[20] = fifoOut[48][2];
              muxOutConnector[21] = fifoOut[49][2];
              muxOutConnector[22] = fifoOut[50][2];
              muxOutConnector[23] = fifoOut[51][2];
              muxOutConnector[24] = fifoOut[26][1];
              muxOutConnector[25] = fifoOut[27][1];
              muxOutConnector[26] = fifoOut[27][6];
              muxOutConnector[27] = fifoOut[28][6];
              muxOutConnector[28] = fifoOut[29][6];
              muxOutConnector[29] = fifoOut[30][6];
              muxOutConnector[30] = fifoOut[31][6];
              muxOutConnector[31] = fifoOut[32][6];
              muxOutConnector[32] = fifoOut[33][6];
              muxOutConnector[33] = fifoOut[34][6];
              muxOutConnector[34] = fifoOut[35][6];
              muxOutConnector[35] = fifoOut[36][6];
              muxOutConnector[36] = fifoOut[37][6];
              muxOutConnector[37] = fifoOut[38][6];
              muxOutConnector[38] = fifoOut[39][6];
              muxOutConnector[39] = fifoOut[40][6];
              muxOutConnector[40] = fifoOut[41][6];
              muxOutConnector[41] = fifoOut[42][6];
              muxOutConnector[42] = fifoOut[43][6];
              muxOutConnector[43] = fifoOut[44][6];
              muxOutConnector[44] = fifoOut[45][6];
              muxOutConnector[45] = fifoOut[46][6];
              muxOutConnector[46] = fifoOut[47][6];
              muxOutConnector[47] = fifoOut[48][6];
              muxOutConnector[48] = fifoOut[49][6];
              muxOutConnector[49] = fifoOut[50][6];
              muxOutConnector[50] = fifoOut[51][6];
              muxOutConnector[51] = fifoOut[26][5];
       end
       4: begin
              muxOutConnector[0] = fifoOut[28][2];
              muxOutConnector[1] = fifoOut[29][2];
              muxOutConnector[2] = fifoOut[30][2];
              muxOutConnector[3] = fifoOut[31][2];
              muxOutConnector[4] = fifoOut[32][2];
              muxOutConnector[5] = fifoOut[33][2];
              muxOutConnector[6] = fifoOut[34][2];
              muxOutConnector[7] = fifoOut[35][2];
              muxOutConnector[8] = fifoOut[36][2];
              muxOutConnector[9] = fifoOut[37][2];
              muxOutConnector[10] = fifoOut[38][2];
              muxOutConnector[11] = fifoOut[39][2];
              muxOutConnector[12] = fifoOut[40][2];
              muxOutConnector[13] = fifoOut[41][2];
              muxOutConnector[14] = fifoOut[42][2];
              muxOutConnector[15] = fifoOut[43][2];
              muxOutConnector[16] = fifoOut[44][2];
              muxOutConnector[17] = fifoOut[45][2];
              muxOutConnector[18] = fifoOut[46][2];
              muxOutConnector[19] = fifoOut[47][2];
              muxOutConnector[20] = fifoOut[48][2];
              muxOutConnector[21] = fifoOut[49][2];
              muxOutConnector[22] = fifoOut[50][2];
              muxOutConnector[23] = fifoOut[51][2];
              muxOutConnector[24] = fifoOut[26][1];
              muxOutConnector[25] = fifoOut[27][1];
              muxOutConnector[26] = fifoOut[27][6];
              muxOutConnector[27] = fifoOut[28][6];
              muxOutConnector[28] = fifoOut[29][6];
              muxOutConnector[29] = fifoOut[30][6];
              muxOutConnector[30] = fifoOut[31][6];
              muxOutConnector[31] = fifoOut[32][6];
              muxOutConnector[32] = fifoOut[33][6];
              muxOutConnector[33] = fifoOut[34][6];
              muxOutConnector[34] = fifoOut[35][6];
              muxOutConnector[35] = fifoOut[36][6];
              muxOutConnector[36] = fifoOut[37][6];
              muxOutConnector[37] = fifoOut[38][6];
              muxOutConnector[38] = fifoOut[39][6];
              muxOutConnector[39] = fifoOut[40][6];
              muxOutConnector[40] = fifoOut[41][6];
              muxOutConnector[41] = fifoOut[42][6];
              muxOutConnector[42] = fifoOut[43][6];
              muxOutConnector[43] = fifoOut[44][6];
              muxOutConnector[44] = fifoOut[45][6];
              muxOutConnector[45] = fifoOut[46][6];
              muxOutConnector[46] = fifoOut[47][6];
              muxOutConnector[47] = fifoOut[48][6];
              muxOutConnector[48] = fifoOut[49][6];
              muxOutConnector[49] = fifoOut[50][6];
              muxOutConnector[50] = fifoOut[51][6];
              muxOutConnector[51] = fifoOut[26][5];
       end
       5: begin
              muxOutConnector[0] = fifoOut[28][2];
              muxOutConnector[1] = fifoOut[29][2];
              muxOutConnector[2] = fifoOut[30][2];
              muxOutConnector[3] = fifoOut[31][2];
              muxOutConnector[4] = fifoOut[32][2];
              muxOutConnector[5] = fifoOut[33][2];
              muxOutConnector[6] = fifoOut[34][2];
              muxOutConnector[7] = fifoOut[35][2];
              muxOutConnector[8] = fifoOut[36][2];
              muxOutConnector[9] = fifoOut[37][2];
              muxOutConnector[10] = fifoOut[38][2];
              muxOutConnector[11] = fifoOut[39][2];
              muxOutConnector[12] = fifoOut[40][2];
              muxOutConnector[13] = fifoOut[41][2];
              muxOutConnector[14] = fifoOut[42][2];
              muxOutConnector[15] = fifoOut[43][2];
              muxOutConnector[16] = fifoOut[44][2];
              muxOutConnector[17] = fifoOut[45][2];
              muxOutConnector[18] = fifoOut[46][2];
              muxOutConnector[19] = fifoOut[47][2];
              muxOutConnector[20] = fifoOut[48][2];
              muxOutConnector[21] = fifoOut[49][2];
              muxOutConnector[22] = fifoOut[50][2];
              muxOutConnector[23] = fifoOut[51][2];
              muxOutConnector[24] = fifoOut[26][1];
              muxOutConnector[25] = fifoOut[27][1];
              muxOutConnector[26] = fifoOut[27][6];
              muxOutConnector[27] = fifoOut[28][6];
              muxOutConnector[28] = fifoOut[29][6];
              muxOutConnector[29] = fifoOut[30][6];
              muxOutConnector[30] = fifoOut[31][6];
              muxOutConnector[31] = fifoOut[32][6];
              muxOutConnector[32] = fifoOut[33][6];
              muxOutConnector[33] = fifoOut[34][6];
              muxOutConnector[34] = fifoOut[35][6];
              muxOutConnector[35] = fifoOut[36][6];
              muxOutConnector[36] = fifoOut[37][6];
              muxOutConnector[37] = fifoOut[38][6];
              muxOutConnector[38] = fifoOut[39][6];
              muxOutConnector[39] = fifoOut[40][6];
              muxOutConnector[40] = fifoOut[41][6];
              muxOutConnector[41] = fifoOut[42][6];
              muxOutConnector[42] = fifoOut[43][6];
              muxOutConnector[43] = fifoOut[44][6];
              muxOutConnector[44] = fifoOut[45][6];
              muxOutConnector[45] = fifoOut[46][6];
              muxOutConnector[46] = fifoOut[47][6];
              muxOutConnector[47] = fifoOut[48][6];
              muxOutConnector[48] = fifoOut[49][6];
              muxOutConnector[49] = fifoOut[50][6];
              muxOutConnector[50] = fifoOut[51][6];
              muxOutConnector[51] = fifoOut[26][5];
       end
       6: begin
              muxOutConnector[0] = fifoOut[28][2];
              muxOutConnector[1] = fifoOut[29][2];
              muxOutConnector[2] = fifoOut[30][2];
              muxOutConnector[3] = fifoOut[31][2];
              muxOutConnector[4] = fifoOut[32][2];
              muxOutConnector[5] = fifoOut[33][2];
              muxOutConnector[6] = fifoOut[34][2];
              muxOutConnector[7] = fifoOut[35][2];
              muxOutConnector[8] = fifoOut[36][2];
              muxOutConnector[9] = fifoOut[37][2];
              muxOutConnector[10] = fifoOut[38][2];
              muxOutConnector[11] = fifoOut[39][2];
              muxOutConnector[12] = fifoOut[40][2];
              muxOutConnector[13] = fifoOut[41][2];
              muxOutConnector[14] = fifoOut[42][2];
              muxOutConnector[15] = fifoOut[43][2];
              muxOutConnector[16] = fifoOut[44][2];
              muxOutConnector[17] = fifoOut[45][2];
              muxOutConnector[18] = fifoOut[46][2];
              muxOutConnector[19] = fifoOut[47][2];
              muxOutConnector[20] = fifoOut[48][2];
              muxOutConnector[21] = fifoOut[49][2];
              muxOutConnector[22] = fifoOut[50][2];
              muxOutConnector[23] = fifoOut[51][2];
              muxOutConnector[24] = fifoOut[26][1];
              muxOutConnector[25] = fifoOut[27][1];
              muxOutConnector[26] = fifoOut[27][6];
              muxOutConnector[27] = fifoOut[28][6];
              muxOutConnector[28] = fifoOut[29][6];
              muxOutConnector[29] = fifoOut[30][6];
              muxOutConnector[30] = fifoOut[31][6];
              muxOutConnector[31] = fifoOut[32][6];
              muxOutConnector[32] = fifoOut[33][6];
              muxOutConnector[33] = fifoOut[34][6];
              muxOutConnector[34] = fifoOut[35][6];
              muxOutConnector[35] = fifoOut[36][6];
              muxOutConnector[36] = fifoOut[37][6];
              muxOutConnector[37] = fifoOut[38][6];
              muxOutConnector[38] = fifoOut[39][6];
              muxOutConnector[39] = fifoOut[40][6];
              muxOutConnector[40] = fifoOut[41][6];
              muxOutConnector[41] = fifoOut[42][6];
              muxOutConnector[42] = fifoOut[23][3];
              muxOutConnector[43] = fifoOut[24][3];
              muxOutConnector[44] = fifoOut[25][3];
              muxOutConnector[45] = fifoOut[0][2];
              muxOutConnector[46] = fifoOut[1][2];
              muxOutConnector[47] = fifoOut[2][2];
              muxOutConnector[48] = fifoOut[3][2];
              muxOutConnector[49] = fifoOut[4][2];
              muxOutConnector[50] = fifoOut[5][2];
              muxOutConnector[51] = fifoOut[6][2];
       end
       7: begin
              muxOutConnector[0] = fifoOut[28][2];
              muxOutConnector[1] = fifoOut[29][2];
              muxOutConnector[2] = fifoOut[30][2];
              muxOutConnector[3] = fifoOut[31][2];
              muxOutConnector[4] = fifoOut[32][2];
              muxOutConnector[5] = fifoOut[33][2];
              muxOutConnector[6] = fifoOut[34][2];
              muxOutConnector[7] = fifoOut[35][2];
              muxOutConnector[8] = fifoOut[36][2];
              muxOutConnector[9] = fifoOut[37][2];
              muxOutConnector[10] = fifoOut[38][2];
              muxOutConnector[11] = fifoOut[39][2];
              muxOutConnector[12] = fifoOut[40][2];
              muxOutConnector[13] = fifoOut[41][2];
              muxOutConnector[14] = fifoOut[42][2];
              muxOutConnector[15] = fifoOut[43][2];
              muxOutConnector[16] = fifoOut[44][2];
              muxOutConnector[17] = fifoOut[45][2];
              muxOutConnector[18] = fifoOut[46][2];
              muxOutConnector[19] = fifoOut[47][2];
              muxOutConnector[20] = fifoOut[48][2];
              muxOutConnector[21] = fifoOut[49][2];
              muxOutConnector[22] = fifoOut[50][2];
              muxOutConnector[23] = fifoOut[51][2];
              muxOutConnector[24] = fifoOut[26][1];
              muxOutConnector[25] = fifoOut[27][1];
              muxOutConnector[26] = fifoOut[7][3];
              muxOutConnector[27] = fifoOut[8][3];
              muxOutConnector[28] = fifoOut[9][3];
              muxOutConnector[29] = fifoOut[10][3];
              muxOutConnector[30] = fifoOut[11][3];
              muxOutConnector[31] = fifoOut[12][3];
              muxOutConnector[32] = fifoOut[13][3];
              muxOutConnector[33] = fifoOut[14][3];
              muxOutConnector[34] = fifoOut[15][3];
              muxOutConnector[35] = fifoOut[16][3];
              muxOutConnector[36] = fifoOut[17][3];
              muxOutConnector[37] = fifoOut[18][3];
              muxOutConnector[38] = fifoOut[19][3];
              muxOutConnector[39] = fifoOut[20][3];
              muxOutConnector[40] = fifoOut[21][3];
              muxOutConnector[41] = fifoOut[22][3];
              muxOutConnector[42] = fifoOut[23][3];
              muxOutConnector[43] = fifoOut[24][3];
              muxOutConnector[44] = fifoOut[25][3];
              muxOutConnector[45] = fifoOut[0][2];
              muxOutConnector[46] = fifoOut[1][2];
              muxOutConnector[47] = fifoOut[2][2];
              muxOutConnector[48] = fifoOut[3][2];
              muxOutConnector[49] = fifoOut[4][2];
              muxOutConnector[50] = fifoOut[5][2];
              muxOutConnector[51] = fifoOut[6][2];
       end
       8: begin
              muxOutConnector[0] = fifoOut[28][2];
              muxOutConnector[1] = fifoOut[29][2];
              muxOutConnector[2] = fifoOut[30][2];
              muxOutConnector[3] = fifoOut[31][2];
              muxOutConnector[4] = fifoOut[32][2];
              muxOutConnector[5] = fifoOut[33][2];
              muxOutConnector[6] = fifoOut[34][2];
              muxOutConnector[7] = fifoOut[35][2];
              muxOutConnector[8] = fifoOut[36][2];
              muxOutConnector[9] = fifoOut[37][2];
              muxOutConnector[10] = fifoOut[38][2];
              muxOutConnector[11] = fifoOut[39][2];
              muxOutConnector[12] = fifoOut[40][2];
              muxOutConnector[13] = fifoOut[41][2];
              muxOutConnector[14] = fifoOut[42][2];
              muxOutConnector[15] = fifoOut[43][2];
              muxOutConnector[16] = fifoOut[44][2];
              muxOutConnector[17] = fifoOut[45][2];
              muxOutConnector[18] = fifoOut[46][2];
              muxOutConnector[19] = fifoOut[47][2];
              muxOutConnector[20] = fifoOut[48][2];
              muxOutConnector[21] = fifoOut[49][2];
              muxOutConnector[22] = fifoOut[50][2];
              muxOutConnector[23] = fifoOut[51][2];
              muxOutConnector[24] = fifoOut[26][1];
              muxOutConnector[25] = fifoOut[27][1];
              muxOutConnector[26] = fifoOut[7][3];
              muxOutConnector[27] = fifoOut[8][3];
              muxOutConnector[28] = fifoOut[9][3];
              muxOutConnector[29] = fifoOut[10][3];
              muxOutConnector[30] = fifoOut[11][3];
              muxOutConnector[31] = fifoOut[12][3];
              muxOutConnector[32] = fifoOut[13][3];
              muxOutConnector[33] = fifoOut[14][3];
              muxOutConnector[34] = fifoOut[15][3];
              muxOutConnector[35] = fifoOut[16][3];
              muxOutConnector[36] = fifoOut[17][3];
              muxOutConnector[37] = fifoOut[18][3];
              muxOutConnector[38] = fifoOut[19][3];
              muxOutConnector[39] = fifoOut[20][3];
              muxOutConnector[40] = fifoOut[21][3];
              muxOutConnector[41] = fifoOut[22][3];
              muxOutConnector[42] = fifoOut[23][3];
              muxOutConnector[43] = fifoOut[24][3];
              muxOutConnector[44] = fifoOut[25][3];
              muxOutConnector[45] = fifoOut[0][2];
              muxOutConnector[46] = fifoOut[1][2];
              muxOutConnector[47] = fifoOut[2][2];
              muxOutConnector[48] = fifoOut[3][2];
              muxOutConnector[49] = fifoOut[4][2];
              muxOutConnector[50] = fifoOut[5][2];
              muxOutConnector[51] = fifoOut[6][2];
       end
       9: begin
              muxOutConnector[0] = fifoOut[28][2];
              muxOutConnector[1] = fifoOut[29][2];
              muxOutConnector[2] = fifoOut[30][2];
              muxOutConnector[3] = fifoOut[31][2];
              muxOutConnector[4] = fifoOut[32][2];
              muxOutConnector[5] = fifoOut[33][2];
              muxOutConnector[6] = fifoOut[34][2];
              muxOutConnector[7] = fifoOut[35][2];
              muxOutConnector[8] = fifoOut[36][2];
              muxOutConnector[9] = fifoOut[37][2];
              muxOutConnector[10] = fifoOut[38][2];
              muxOutConnector[11] = fifoOut[39][2];
              muxOutConnector[12] = fifoOut[40][2];
              muxOutConnector[13] = fifoOut[41][2];
              muxOutConnector[14] = fifoOut[42][2];
              muxOutConnector[15] = fifoOut[43][2];
              muxOutConnector[16] = fifoOut[44][2];
              muxOutConnector[17] = fifoOut[45][2];
              muxOutConnector[18] = fifoOut[46][2];
              muxOutConnector[19] = fifoOut[47][2];
              muxOutConnector[20] = fifoOut[48][2];
              muxOutConnector[21] = fifoOut[49][2];
              muxOutConnector[22] = fifoOut[50][2];
              muxOutConnector[23] = fifoOut[51][2];
              muxOutConnector[24] = fifoOut[26][1];
              muxOutConnector[25] = fifoOut[27][1];
              muxOutConnector[26] = fifoOut[7][3];
              muxOutConnector[27] = fifoOut[8][3];
              muxOutConnector[28] = fifoOut[9][3];
              muxOutConnector[29] = fifoOut[10][3];
              muxOutConnector[30] = fifoOut[11][3];
              muxOutConnector[31] = fifoOut[12][3];
              muxOutConnector[32] = fifoOut[13][3];
              muxOutConnector[33] = fifoOut[14][3];
              muxOutConnector[34] = fifoOut[15][3];
              muxOutConnector[35] = fifoOut[16][3];
              muxOutConnector[36] = fifoOut[17][3];
              muxOutConnector[37] = fifoOut[18][3];
              muxOutConnector[38] = fifoOut[19][3];
              muxOutConnector[39] = fifoOut[20][3];
              muxOutConnector[40] = fifoOut[21][3];
              muxOutConnector[41] = fifoOut[22][3];
              muxOutConnector[42] = fifoOut[23][3];
              muxOutConnector[43] = fifoOut[24][3];
              muxOutConnector[44] = fifoOut[25][3];
              muxOutConnector[45] = fifoOut[0][2];
              muxOutConnector[46] = fifoOut[1][2];
              muxOutConnector[47] = fifoOut[2][2];
              muxOutConnector[48] = fifoOut[3][2];
              muxOutConnector[49] = fifoOut[4][2];
              muxOutConnector[50] = fifoOut[5][2];
              muxOutConnector[51] = fifoOut[6][2];
       end
       10: begin
              muxOutConnector[0] = fifoOut[28][2];
              muxOutConnector[1] = fifoOut[29][2];
              muxOutConnector[2] = fifoOut[30][2];
              muxOutConnector[3] = fifoOut[31][2];
              muxOutConnector[4] = fifoOut[32][2];
              muxOutConnector[5] = fifoOut[33][2];
              muxOutConnector[6] = fifoOut[34][2];
              muxOutConnector[7] = fifoOut[35][2];
              muxOutConnector[8] = fifoOut[36][2];
              muxOutConnector[9] = fifoOut[37][2];
              muxOutConnector[10] = fifoOut[38][2];
              muxOutConnector[11] = fifoOut[39][2];
              muxOutConnector[12] = fifoOut[40][2];
              muxOutConnector[13] = fifoOut[41][2];
              muxOutConnector[14] = fifoOut[42][2];
              muxOutConnector[15] = fifoOut[43][2];
              muxOutConnector[16] = fifoOut[44][2];
              muxOutConnector[17] = fifoOut[45][2];
              muxOutConnector[18] = fifoOut[46][2];
              muxOutConnector[19] = fifoOut[47][2];
              muxOutConnector[20] = fifoOut[48][2];
              muxOutConnector[21] = fifoOut[49][2];
              muxOutConnector[22] = fifoOut[50][2];
              muxOutConnector[23] = fifoOut[51][2];
              muxOutConnector[24] = fifoOut[26][1];
              muxOutConnector[25] = fifoOut[27][1];
              muxOutConnector[26] = fifoOut[7][3];
              muxOutConnector[27] = fifoOut[8][3];
              muxOutConnector[28] = fifoOut[9][3];
              muxOutConnector[29] = fifoOut[10][3];
              muxOutConnector[30] = fifoOut[11][3];
              muxOutConnector[31] = fifoOut[12][3];
              muxOutConnector[32] = fifoOut[13][3];
              muxOutConnector[33] = fifoOut[14][3];
              muxOutConnector[34] = fifoOut[15][3];
              muxOutConnector[35] = fifoOut[16][3];
              muxOutConnector[36] = fifoOut[17][3];
              muxOutConnector[37] = fifoOut[18][3];
              muxOutConnector[38] = fifoOut[19][3];
              muxOutConnector[39] = fifoOut[20][3];
              muxOutConnector[40] = fifoOut[21][3];
              muxOutConnector[41] = fifoOut[22][3];
              muxOutConnector[42] = fifoOut[23][3];
              muxOutConnector[43] = fifoOut[24][3];
              muxOutConnector[44] = fifoOut[25][3];
              muxOutConnector[45] = fifoOut[0][2];
              muxOutConnector[46] = fifoOut[1][2];
              muxOutConnector[47] = fifoOut[2][2];
              muxOutConnector[48] = fifoOut[3][2];
              muxOutConnector[49] = fifoOut[4][2];
              muxOutConnector[50] = fifoOut[5][2];
              muxOutConnector[51] = fifoOut[6][2];
       end
       11: begin
              muxOutConnector[0] = fifoOut[28][2];
              muxOutConnector[1] = fifoOut[29][2];
              muxOutConnector[2] = fifoOut[30][2];
              muxOutConnector[3] = fifoOut[31][2];
              muxOutConnector[4] = fifoOut[32][2];
              muxOutConnector[5] = fifoOut[33][2];
              muxOutConnector[6] = fifoOut[34][2];
              muxOutConnector[7] = fifoOut[35][2];
              muxOutConnector[8] = fifoOut[36][2];
              muxOutConnector[9] = fifoOut[37][2];
              muxOutConnector[10] = fifoOut[38][2];
              muxOutConnector[11] = fifoOut[39][2];
              muxOutConnector[12] = fifoOut[40][2];
              muxOutConnector[13] = fifoOut[41][2];
              muxOutConnector[14] = fifoOut[42][2];
              muxOutConnector[15] = fifoOut[43][2];
              muxOutConnector[16] = fifoOut[44][2];
              muxOutConnector[17] = fifoOut[45][2];
              muxOutConnector[18] = fifoOut[0][10];
              muxOutConnector[19] = fifoOut[1][10];
              muxOutConnector[20] = fifoOut[2][10];
              muxOutConnector[21] = fifoOut[3][10];
              muxOutConnector[22] = fifoOut[4][10];
              muxOutConnector[23] = fifoOut[5][10];
              muxOutConnector[24] = fifoOut[6][10];
              muxOutConnector[25] = fifoOut[7][10];
              muxOutConnector[26] = fifoOut[7][3];
              muxOutConnector[27] = fifoOut[8][3];
              muxOutConnector[28] = fifoOut[9][3];
              muxOutConnector[29] = fifoOut[10][3];
              muxOutConnector[30] = fifoOut[11][3];
              muxOutConnector[31] = fifoOut[12][3];
              muxOutConnector[32] = fifoOut[13][3];
              muxOutConnector[33] = fifoOut[14][3];
              muxOutConnector[34] = fifoOut[15][3];
              muxOutConnector[35] = fifoOut[16][3];
              muxOutConnector[36] = fifoOut[17][3];
              muxOutConnector[37] = fifoOut[18][3];
              muxOutConnector[38] = fifoOut[19][3];
              muxOutConnector[39] = fifoOut[20][3];
              muxOutConnector[40] = fifoOut[21][3];
              muxOutConnector[41] = fifoOut[22][3];
              muxOutConnector[42] = fifoOut[23][3];
              muxOutConnector[43] = fifoOut[24][3];
              muxOutConnector[44] = fifoOut[25][3];
              muxOutConnector[45] = fifoOut[0][2];
              muxOutConnector[46] = fifoOut[1][2];
              muxOutConnector[47] = fifoOut[2][2];
              muxOutConnector[48] = fifoOut[3][2];
              muxOutConnector[49] = fifoOut[4][2];
              muxOutConnector[50] = fifoOut[5][2];
              muxOutConnector[51] = fifoOut[6][2];
       end
       12: begin
              muxOutConnector[0] = fifoOut[8][11];
              muxOutConnector[1] = fifoOut[9][11];
              muxOutConnector[2] = fifoOut[10][11];
              muxOutConnector[3] = fifoOut[11][11];
              muxOutConnector[4] = fifoOut[12][11];
              muxOutConnector[5] = fifoOut[13][11];
              muxOutConnector[6] = fifoOut[14][11];
              muxOutConnector[7] = fifoOut[15][11];
              muxOutConnector[8] = fifoOut[16][11];
              muxOutConnector[9] = fifoOut[17][11];
              muxOutConnector[10] = fifoOut[18][11];
              muxOutConnector[11] = fifoOut[19][11];
              muxOutConnector[12] = fifoOut[20][11];
              muxOutConnector[13] = fifoOut[21][11];
              muxOutConnector[14] = fifoOut[22][11];
              muxOutConnector[15] = fifoOut[23][11];
              muxOutConnector[16] = fifoOut[24][11];
              muxOutConnector[17] = fifoOut[25][11];
              muxOutConnector[18] = fifoOut[0][10];
              muxOutConnector[19] = fifoOut[1][10];
              muxOutConnector[20] = fifoOut[2][10];
              muxOutConnector[21] = fifoOut[3][10];
              muxOutConnector[22] = fifoOut[4][10];
              muxOutConnector[23] = fifoOut[5][10];
              muxOutConnector[24] = fifoOut[6][10];
              muxOutConnector[25] = fifoOut[7][10];
              muxOutConnector[26] = fifoOut[7][3];
              muxOutConnector[27] = fifoOut[8][3];
              muxOutConnector[28] = fifoOut[9][3];
              muxOutConnector[29] = fifoOut[10][3];
              muxOutConnector[30] = fifoOut[11][3];
              muxOutConnector[31] = fifoOut[12][3];
              muxOutConnector[32] = fifoOut[13][3];
              muxOutConnector[33] = fifoOut[14][3];
              muxOutConnector[34] = fifoOut[15][3];
              muxOutConnector[35] = fifoOut[16][3];
              muxOutConnector[36] = fifoOut[17][3];
              muxOutConnector[37] = fifoOut[18][3];
              muxOutConnector[38] = fifoOut[19][3];
              muxOutConnector[39] = fifoOut[20][3];
              muxOutConnector[40] = fifoOut[21][3];
              muxOutConnector[41] = fifoOut[22][3];
              muxOutConnector[42] = fifoOut[23][3];
              muxOutConnector[43] = fifoOut[24][3];
              muxOutConnector[44] = fifoOut[25][3];
              muxOutConnector[45] = fifoOut[0][2];
              muxOutConnector[46] = fifoOut[1][2];
              muxOutConnector[47] = fifoOut[2][2];
              muxOutConnector[48] = fifoOut[3][2];
              muxOutConnector[49] = fifoOut[4][2];
              muxOutConnector[50] = fifoOut[5][2];
              muxOutConnector[51] = fifoOut[6][2];
       end
       13: begin
              muxOutConnector[0] = fifoOut[8][11];
              muxOutConnector[1] = fifoOut[9][11];
              muxOutConnector[2] = fifoOut[10][11];
              muxOutConnector[3] = fifoOut[11][11];
              muxOutConnector[4] = fifoOut[12][11];
              muxOutConnector[5] = fifoOut[13][11];
              muxOutConnector[6] = fifoOut[14][11];
              muxOutConnector[7] = fifoOut[15][11];
              muxOutConnector[8] = fifoOut[16][11];
              muxOutConnector[9] = fifoOut[17][11];
              muxOutConnector[10] = fifoOut[18][11];
              muxOutConnector[11] = fifoOut[19][11];
              muxOutConnector[12] = fifoOut[20][11];
              muxOutConnector[13] = fifoOut[21][11];
              muxOutConnector[14] = fifoOut[22][11];
              muxOutConnector[15] = fifoOut[23][11];
              muxOutConnector[16] = fifoOut[24][11];
              muxOutConnector[17] = fifoOut[25][11];
              muxOutConnector[18] = fifoOut[0][10];
              muxOutConnector[19] = fifoOut[1][10];
              muxOutConnector[20] = fifoOut[2][10];
              muxOutConnector[21] = fifoOut[3][10];
              muxOutConnector[22] = fifoOut[4][10];
              muxOutConnector[23] = fifoOut[5][10];
              muxOutConnector[24] = fifoOut[6][10];
              muxOutConnector[25] = fifoOut[7][10];
              muxOutConnector[26] = fifoOut[7][3];
              muxOutConnector[27] = fifoOut[8][3];
              muxOutConnector[28] = fifoOut[9][3];
              muxOutConnector[29] = fifoOut[10][3];
              muxOutConnector[30] = fifoOut[11][3];
              muxOutConnector[31] = fifoOut[12][3];
              muxOutConnector[32] = fifoOut[13][3];
              muxOutConnector[33] = fifoOut[14][3];
              muxOutConnector[34] = fifoOut[15][3];
              muxOutConnector[35] = fifoOut[16][3];
              muxOutConnector[36] = fifoOut[17][3];
              muxOutConnector[37] = fifoOut[18][3];
              muxOutConnector[38] = fifoOut[19][3];
              muxOutConnector[39] = fifoOut[20][3];
              muxOutConnector[40] = fifoOut[21][3];
              muxOutConnector[41] = fifoOut[22][3];
              muxOutConnector[42] = fifoOut[23][3];
              muxOutConnector[43] = fifoOut[24][3];
              muxOutConnector[44] = fifoOut[25][3];
              muxOutConnector[45] = fifoOut[0][2];
              muxOutConnector[46] = fifoOut[1][2];
              muxOutConnector[47] = fifoOut[2][2];
              muxOutConnector[48] = fifoOut[3][2];
              muxOutConnector[49] = fifoOut[4][2];
              muxOutConnector[50] = fifoOut[5][2];
              muxOutConnector[51] = fifoOut[6][2];
       end
       14: begin
              muxOutConnector[0] = fifoOut[8][11];
              muxOutConnector[1] = fifoOut[9][11];
              muxOutConnector[2] = fifoOut[10][11];
              muxOutConnector[3] = fifoOut[11][11];
              muxOutConnector[4] = fifoOut[12][11];
              muxOutConnector[5] = fifoOut[13][11];
              muxOutConnector[6] = fifoOut[14][11];
              muxOutConnector[7] = fifoOut[15][11];
              muxOutConnector[8] = fifoOut[16][11];
              muxOutConnector[9] = fifoOut[17][11];
              muxOutConnector[10] = fifoOut[18][11];
              muxOutConnector[11] = fifoOut[19][11];
              muxOutConnector[12] = fifoOut[20][11];
              muxOutConnector[13] = fifoOut[21][11];
              muxOutConnector[14] = fifoOut[22][11];
              muxOutConnector[15] = fifoOut[23][11];
              muxOutConnector[16] = fifoOut[24][11];
              muxOutConnector[17] = fifoOut[25][11];
              muxOutConnector[18] = fifoOut[0][10];
              muxOutConnector[19] = fifoOut[1][10];
              muxOutConnector[20] = fifoOut[2][10];
              muxOutConnector[21] = fifoOut[3][10];
              muxOutConnector[22] = fifoOut[4][10];
              muxOutConnector[23] = fifoOut[5][10];
              muxOutConnector[24] = fifoOut[6][10];
              muxOutConnector[25] = fifoOut[7][10];
              muxOutConnector[26] = fifoOut[7][3];
              muxOutConnector[27] = fifoOut[8][3];
              muxOutConnector[28] = fifoOut[9][3];
              muxOutConnector[29] = fifoOut[10][3];
              muxOutConnector[30] = fifoOut[11][3];
              muxOutConnector[31] = fifoOut[12][3];
              muxOutConnector[32] = fifoOut[13][3];
              muxOutConnector[33] = fifoOut[14][3];
              muxOutConnector[34] = fifoOut[15][3];
              muxOutConnector[35] = fifoOut[16][3];
              muxOutConnector[36] = fifoOut[17][3];
              muxOutConnector[37] = fifoOut[18][3];
              muxOutConnector[38] = fifoOut[19][3];
              muxOutConnector[39] = fifoOut[20][3];
              muxOutConnector[40] = fifoOut[21][3];
              muxOutConnector[41] = fifoOut[22][3];
              muxOutConnector[42] = fifoOut[23][3];
              muxOutConnector[43] = fifoOut[24][3];
              muxOutConnector[44] = fifoOut[25][3];
              muxOutConnector[45] = fifoOut[0][2];
              muxOutConnector[46] = fifoOut[1][2];
              muxOutConnector[47] = fifoOut[2][2];
              muxOutConnector[48] = fifoOut[3][2];
              muxOutConnector[49] = fifoOut[4][2];
              muxOutConnector[50] = fifoOut[5][2];
              muxOutConnector[51] = fifoOut[6][2];
       end
       15: begin
              muxOutConnector[0] = fifoOut[8][11];
              muxOutConnector[1] = fifoOut[9][11];
              muxOutConnector[2] = fifoOut[10][11];
              muxOutConnector[3] = fifoOut[11][11];
              muxOutConnector[4] = fifoOut[12][11];
              muxOutConnector[5] = fifoOut[13][11];
              muxOutConnector[6] = fifoOut[14][11];
              muxOutConnector[7] = fifoOut[15][11];
              muxOutConnector[8] = fifoOut[16][11];
              muxOutConnector[9] = fifoOut[17][11];
              muxOutConnector[10] = fifoOut[18][11];
              muxOutConnector[11] = fifoOut[19][11];
              muxOutConnector[12] = fifoOut[20][11];
              muxOutConnector[13] = fifoOut[21][11];
              muxOutConnector[14] = fifoOut[22][11];
              muxOutConnector[15] = fifoOut[23][11];
              muxOutConnector[16] = fifoOut[24][11];
              muxOutConnector[17] = fifoOut[25][11];
              muxOutConnector[18] = fifoOut[0][10];
              muxOutConnector[19] = fifoOut[1][10];
              muxOutConnector[20] = fifoOut[2][10];
              muxOutConnector[21] = fifoOut[3][10];
              muxOutConnector[22] = fifoOut[4][10];
              muxOutConnector[23] = fifoOut[5][10];
              muxOutConnector[24] = fifoOut[6][10];
              muxOutConnector[25] = fifoOut[7][10];
              muxOutConnector[26] = fifoOut[7][3];
              muxOutConnector[27] = fifoOut[8][3];
              muxOutConnector[28] = fifoOut[9][3];
              muxOutConnector[29] = fifoOut[10][3];
              muxOutConnector[30] = fifoOut[11][3];
              muxOutConnector[31] = fifoOut[12][3];
              muxOutConnector[32] = fifoOut[13][3];
              muxOutConnector[33] = fifoOut[14][3];
              muxOutConnector[34] = fifoOut[15][3];
              muxOutConnector[35] = fifoOut[16][3];
              muxOutConnector[36] = fifoOut[46][2];
              muxOutConnector[37] = fifoOut[47][2];
              muxOutConnector[38] = fifoOut[48][2];
              muxOutConnector[39] = fifoOut[49][2];
              muxOutConnector[40] = fifoOut[50][2];
              muxOutConnector[41] = fifoOut[51][2];
              muxOutConnector[42] = fifoOut[26][1];
              muxOutConnector[43] = fifoOut[27][1];
              muxOutConnector[44] = fifoOut[28][1];
              muxOutConnector[45] = fifoOut[29][1];
              muxOutConnector[46] = fifoOut[30][1];
              muxOutConnector[47] = fifoOut[31][1];
              muxOutConnector[48] = fifoOut[32][1];
              muxOutConnector[49] = fifoOut[33][1];
              muxOutConnector[50] = fifoOut[34][1];
              muxOutConnector[51] = fifoOut[35][1];
       end
       16: begin
              muxOutConnector[0] = fifoOut[8][11];
              muxOutConnector[1] = fifoOut[9][11];
              muxOutConnector[2] = fifoOut[10][11];
              muxOutConnector[3] = fifoOut[11][11];
              muxOutConnector[4] = fifoOut[12][11];
              muxOutConnector[5] = fifoOut[13][11];
              muxOutConnector[6] = fifoOut[14][11];
              muxOutConnector[7] = fifoOut[15][11];
              muxOutConnector[8] = fifoOut[16][11];
              muxOutConnector[9] = fifoOut[17][11];
              muxOutConnector[10] = fifoOut[18][11];
              muxOutConnector[11] = fifoOut[19][11];
              muxOutConnector[12] = fifoOut[20][11];
              muxOutConnector[13] = fifoOut[21][11];
              muxOutConnector[14] = fifoOut[22][11];
              muxOutConnector[15] = fifoOut[23][11];
              muxOutConnector[16] = fifoOut[24][11];
              muxOutConnector[17] = fifoOut[25][11];
              muxOutConnector[18] = fifoOut[0][10];
              muxOutConnector[19] = fifoOut[1][10];
              muxOutConnector[20] = fifoOut[2][10];
              muxOutConnector[21] = fifoOut[3][10];
              muxOutConnector[22] = fifoOut[4][10];
              muxOutConnector[23] = fifoOut[5][10];
              muxOutConnector[24] = fifoOut[6][10];
              muxOutConnector[25] = fifoOut[7][10];
              muxOutConnector[26] = fifoOut[36][2];
              muxOutConnector[27] = fifoOut[37][2];
              muxOutConnector[28] = fifoOut[38][2];
              muxOutConnector[29] = fifoOut[39][2];
              muxOutConnector[30] = fifoOut[40][2];
              muxOutConnector[31] = fifoOut[41][2];
              muxOutConnector[32] = fifoOut[42][2];
              muxOutConnector[33] = fifoOut[43][2];
              muxOutConnector[34] = fifoOut[44][2];
              muxOutConnector[35] = fifoOut[45][2];
              muxOutConnector[36] = fifoOut[46][2];
              muxOutConnector[37] = fifoOut[47][2];
              muxOutConnector[38] = fifoOut[48][2];
              muxOutConnector[39] = fifoOut[49][2];
              muxOutConnector[40] = fifoOut[50][2];
              muxOutConnector[41] = fifoOut[51][2];
              muxOutConnector[42] = fifoOut[26][1];
              muxOutConnector[43] = fifoOut[27][1];
              muxOutConnector[44] = fifoOut[28][1];
              muxOutConnector[45] = fifoOut[29][1];
              muxOutConnector[46] = fifoOut[30][1];
              muxOutConnector[47] = fifoOut[31][1];
              muxOutConnector[48] = fifoOut[32][1];
              muxOutConnector[49] = fifoOut[33][1];
              muxOutConnector[50] = fifoOut[34][1];
              muxOutConnector[51] = fifoOut[35][1];
       end
       17: begin
              muxOutConnector[0] = fifoOut[8][11];
              muxOutConnector[1] = fifoOut[9][11];
              muxOutConnector[2] = fifoOut[10][11];
              muxOutConnector[3] = fifoOut[11][11];
              muxOutConnector[4] = fifoOut[12][11];
              muxOutConnector[5] = fifoOut[13][11];
              muxOutConnector[6] = fifoOut[14][11];
              muxOutConnector[7] = fifoOut[15][11];
              muxOutConnector[8] = fifoOut[16][11];
              muxOutConnector[9] = fifoOut[17][11];
              muxOutConnector[10] = fifoOut[18][11];
              muxOutConnector[11] = fifoOut[19][11];
              muxOutConnector[12] = fifoOut[20][11];
              muxOutConnector[13] = fifoOut[21][11];
              muxOutConnector[14] = fifoOut[22][11];
              muxOutConnector[15] = fifoOut[23][11];
              muxOutConnector[16] = fifoOut[24][11];
              muxOutConnector[17] = fifoOut[25][11];
              muxOutConnector[18] = fifoOut[0][10];
              muxOutConnector[19] = fifoOut[1][10];
              muxOutConnector[20] = fifoOut[2][10];
              muxOutConnector[21] = fifoOut[3][10];
              muxOutConnector[22] = fifoOut[4][10];
              muxOutConnector[23] = fifoOut[5][10];
              muxOutConnector[24] = fifoOut[6][10];
              muxOutConnector[25] = fifoOut[7][10];
              muxOutConnector[26] = fifoOut[36][2];
              muxOutConnector[27] = fifoOut[37][2];
              muxOutConnector[28] = fifoOut[38][2];
              muxOutConnector[29] = fifoOut[39][2];
              muxOutConnector[30] = fifoOut[40][2];
              muxOutConnector[31] = fifoOut[41][2];
              muxOutConnector[32] = fifoOut[42][2];
              muxOutConnector[33] = fifoOut[43][2];
              muxOutConnector[34] = fifoOut[44][2];
              muxOutConnector[35] = fifoOut[45][2];
              muxOutConnector[36] = fifoOut[46][2];
              muxOutConnector[37] = fifoOut[47][2];
              muxOutConnector[38] = fifoOut[48][2];
              muxOutConnector[39] = fifoOut[49][2];
              muxOutConnector[40] = fifoOut[50][2];
              muxOutConnector[41] = fifoOut[51][2];
              muxOutConnector[42] = fifoOut[26][1];
              muxOutConnector[43] = fifoOut[27][1];
              muxOutConnector[44] = fifoOut[28][1];
              muxOutConnector[45] = fifoOut[29][1];
              muxOutConnector[46] = fifoOut[30][1];
              muxOutConnector[47] = fifoOut[31][1];
              muxOutConnector[48] = fifoOut[32][1];
              muxOutConnector[49] = fifoOut[33][1];
              muxOutConnector[50] = fifoOut[34][1];
              muxOutConnector[51] = fifoOut[35][1];
       end
       18: begin
              muxOutConnector[0] = fifoOut[8][11];
              muxOutConnector[1] = fifoOut[9][11];
              muxOutConnector[2] = fifoOut[10][11];
              muxOutConnector[3] = fifoOut[11][11];
              muxOutConnector[4] = fifoOut[12][11];
              muxOutConnector[5] = fifoOut[13][11];
              muxOutConnector[6] = fifoOut[14][11];
              muxOutConnector[7] = fifoOut[15][11];
              muxOutConnector[8] = fifoOut[16][11];
              muxOutConnector[9] = fifoOut[17][11];
              muxOutConnector[10] = fifoOut[18][11];
              muxOutConnector[11] = fifoOut[19][11];
              muxOutConnector[12] = fifoOut[20][11];
              muxOutConnector[13] = fifoOut[21][11];
              muxOutConnector[14] = fifoOut[22][11];
              muxOutConnector[15] = fifoOut[23][11];
              muxOutConnector[16] = fifoOut[24][11];
              muxOutConnector[17] = fifoOut[25][11];
              muxOutConnector[18] = fifoOut[0][10];
              muxOutConnector[19] = fifoOut[1][10];
              muxOutConnector[20] = fifoOut[2][10];
              muxOutConnector[21] = fifoOut[3][10];
              muxOutConnector[22] = fifoOut[4][10];
              muxOutConnector[23] = fifoOut[5][10];
              muxOutConnector[24] = fifoOut[6][10];
              muxOutConnector[25] = fifoOut[7][10];
              muxOutConnector[26] = fifoOut[36][2];
              muxOutConnector[27] = fifoOut[37][2];
              muxOutConnector[28] = fifoOut[38][2];
              muxOutConnector[29] = fifoOut[39][2];
              muxOutConnector[30] = fifoOut[40][2];
              muxOutConnector[31] = fifoOut[41][2];
              muxOutConnector[32] = fifoOut[42][2];
              muxOutConnector[33] = fifoOut[43][2];
              muxOutConnector[34] = fifoOut[44][2];
              muxOutConnector[35] = fifoOut[45][2];
              muxOutConnector[36] = fifoOut[46][2];
              muxOutConnector[37] = fifoOut[47][2];
              muxOutConnector[38] = fifoOut[48][2];
              muxOutConnector[39] = fifoOut[49][2];
              muxOutConnector[40] = fifoOut[50][2];
              muxOutConnector[41] = fifoOut[51][2];
              muxOutConnector[42] = fifoOut[26][1];
              muxOutConnector[43] = fifoOut[27][1];
              muxOutConnector[44] = fifoOut[28][1];
              muxOutConnector[45] = fifoOut[29][1];
              muxOutConnector[46] = fifoOut[30][1];
              muxOutConnector[47] = fifoOut[31][1];
              muxOutConnector[48] = fifoOut[32][1];
              muxOutConnector[49] = fifoOut[33][1];
              muxOutConnector[50] = fifoOut[34][1];
              muxOutConnector[51] = fifoOut[35][1];
       end
       19: begin
              muxOutConnector[0] = fifoOut[8][11];
              muxOutConnector[1] = fifoOut[9][11];
              muxOutConnector[2] = fifoOut[10][11];
              muxOutConnector[3] = fifoOut[11][11];
              muxOutConnector[4] = fifoOut[12][11];
              muxOutConnector[5] = fifoOut[13][11];
              muxOutConnector[6] = fifoOut[14][11];
              muxOutConnector[7] = fifoOut[15][11];
              muxOutConnector[8] = fifoOut[16][11];
              muxOutConnector[9] = fifoOut[17][11];
              muxOutConnector[10] = fifoOut[18][11];
              muxOutConnector[11] = fifoOut[19][11];
              muxOutConnector[12] = fifoOut[20][11];
              muxOutConnector[13] = fifoOut[21][11];
              muxOutConnector[14] = fifoOut[22][11];
              muxOutConnector[15] = fifoOut[23][11];
              muxOutConnector[16] = fifoOut[24][11];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[36][2];
              muxOutConnector[27] = fifoOut[37][2];
              muxOutConnector[28] = fifoOut[38][2];
              muxOutConnector[29] = fifoOut[39][2];
              muxOutConnector[30] = fifoOut[40][2];
              muxOutConnector[31] = fifoOut[41][2];
              muxOutConnector[32] = fifoOut[42][2];
              muxOutConnector[33] = fifoOut[43][2];
              muxOutConnector[34] = fifoOut[44][2];
              muxOutConnector[35] = fifoOut[45][2];
              muxOutConnector[36] = fifoOut[46][2];
              muxOutConnector[37] = fifoOut[47][2];
              muxOutConnector[38] = fifoOut[48][2];
              muxOutConnector[39] = fifoOut[49][2];
              muxOutConnector[40] = fifoOut[50][2];
              muxOutConnector[41] = fifoOut[51][2];
              muxOutConnector[42] = fifoOut[26][1];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
