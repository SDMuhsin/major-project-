`timescale 1ns / 1ps
module LMem0To1_511_circ14_ys_scripted(
        muxOut,
        ly0In,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 11;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

reg   feedback_en;
reg [ w - 1 : 0 ]column_1[ r - 1 : 0 ];
reg chip_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(chip_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= column_1[i];
         end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
  feedback_en=rd_en;
      if(wr_en)begin
        chip_en=wr_en;
      end
      else begin
        chip_en=feedback_en;
      end
   if(feedback_en)begin
      for(i = r-1; i > -1; i=i-1) begin
        column_1[i] <= fifoOut[i][c-1];
      end
   end
   else begin
      for(i = r-1; i > -1; i=i-1) begin
        column_1[i] <= ly0InConnector[i];
      end
    end
end
always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[29][7];
              muxOutConnector[1] = fifoOut[30][7];
              muxOutConnector[2] = fifoOut[31][7];
              muxOutConnector[3] = fifoOut[32][7];
              muxOutConnector[4] = fifoOut[33][7];
              muxOutConnector[5] = fifoOut[34][7];
              muxOutConnector[6] = fifoOut[35][7];
              muxOutConnector[7] = fifoOut[36][7];
              muxOutConnector[8] = fifoOut[37][7];
              muxOutConnector[9] = fifoOut[38][7];
              muxOutConnector[10] = fifoOut[39][7];
              muxOutConnector[11] = fifoOut[40][7];
              muxOutConnector[12] = fifoOut[41][7];
              muxOutConnector[13] = fifoOut[42][7];
              muxOutConnector[14] = fifoOut[43][7];
              muxOutConnector[15] = fifoOut[44][7];
              muxOutConnector[16] = fifoOut[45][7];
              muxOutConnector[17] = fifoOut[46][7];
              muxOutConnector[18] = fifoOut[47][7];
              muxOutConnector[19] = fifoOut[48][7];
              muxOutConnector[20] = fifoOut[49][7];
              muxOutConnector[21] = fifoOut[50][7];
              muxOutConnector[22] = fifoOut[51][7];
              muxOutConnector[23] = fifoOut[26][6];
              muxOutConnector[24] = fifoOut[27][6];
              muxOutConnector[25] = fifoOut[28][6];
              muxOutConnector[26] = fifoOut[18][5];
              muxOutConnector[27] = fifoOut[19][5];
              muxOutConnector[28] = fifoOut[20][5];
              muxOutConnector[29] = fifoOut[21][5];
              muxOutConnector[30] = fifoOut[22][5];
              muxOutConnector[31] = fifoOut[23][5];
              muxOutConnector[32] = fifoOut[24][5];
              muxOutConnector[33] = fifoOut[25][5];
              muxOutConnector[34] = fifoOut[0][4];
              muxOutConnector[35] = fifoOut[1][4];
              muxOutConnector[36] = fifoOut[2][4];
              muxOutConnector[37] = fifoOut[3][4];
              muxOutConnector[38] = fifoOut[4][4];
              muxOutConnector[39] = fifoOut[5][4];
              muxOutConnector[40] = fifoOut[6][4];
              muxOutConnector[41] = fifoOut[7][4];
              muxOutConnector[42] = fifoOut[8][4];
              muxOutConnector[43] = fifoOut[9][4];
              muxOutConnector[44] = fifoOut[10][4];
              muxOutConnector[45] = fifoOut[11][4];
              muxOutConnector[46] = fifoOut[12][4];
              muxOutConnector[47] = fifoOut[13][4];
              muxOutConnector[48] = fifoOut[14][4];
              muxOutConnector[49] = fifoOut[15][4];
              muxOutConnector[50] = fifoOut[16][4];
              muxOutConnector[51] = fifoOut[17][4];
       end
       1: begin
              muxOutConnector[0] = fifoOut[29][7];
              muxOutConnector[1] = fifoOut[30][7];
              muxOutConnector[2] = fifoOut[31][7];
              muxOutConnector[3] = fifoOut[32][7];
              muxOutConnector[4] = fifoOut[33][7];
              muxOutConnector[5] = fifoOut[34][7];
              muxOutConnector[6] = fifoOut[35][7];
              muxOutConnector[7] = fifoOut[36][7];
              muxOutConnector[8] = fifoOut[37][7];
              muxOutConnector[9] = fifoOut[38][7];
              muxOutConnector[10] = fifoOut[39][7];
              muxOutConnector[11] = fifoOut[40][7];
              muxOutConnector[12] = fifoOut[41][7];
              muxOutConnector[13] = fifoOut[42][7];
              muxOutConnector[14] = fifoOut[43][7];
              muxOutConnector[15] = fifoOut[44][7];
              muxOutConnector[16] = fifoOut[45][7];
              muxOutConnector[17] = fifoOut[46][7];
              muxOutConnector[18] = fifoOut[47][7];
              muxOutConnector[19] = fifoOut[48][7];
              muxOutConnector[20] = fifoOut[49][7];
              muxOutConnector[21] = fifoOut[50][7];
              muxOutConnector[22] = fifoOut[51][7];
              muxOutConnector[23] = fifoOut[26][6];
              muxOutConnector[24] = fifoOut[27][6];
              muxOutConnector[25] = fifoOut[28][6];
              muxOutConnector[26] = fifoOut[18][5];
              muxOutConnector[27] = fifoOut[19][5];
              muxOutConnector[28] = fifoOut[20][5];
              muxOutConnector[29] = fifoOut[21][5];
              muxOutConnector[30] = fifoOut[22][5];
              muxOutConnector[31] = fifoOut[23][5];
              muxOutConnector[32] = fifoOut[24][5];
              muxOutConnector[33] = fifoOut[25][5];
              muxOutConnector[34] = fifoOut[0][4];
              muxOutConnector[35] = fifoOut[1][4];
              muxOutConnector[36] = fifoOut[2][4];
              muxOutConnector[37] = fifoOut[3][4];
              muxOutConnector[38] = fifoOut[4][4];
              muxOutConnector[39] = fifoOut[5][4];
              muxOutConnector[40] = fifoOut[6][4];
              muxOutConnector[41] = fifoOut[7][4];
              muxOutConnector[42] = fifoOut[8][4];
              muxOutConnector[43] = fifoOut[9][4];
              muxOutConnector[44] = fifoOut[10][4];
              muxOutConnector[45] = fifoOut[11][4];
              muxOutConnector[46] = fifoOut[12][4];
              muxOutConnector[47] = fifoOut[13][4];
              muxOutConnector[48] = fifoOut[14][4];
              muxOutConnector[49] = fifoOut[15][4];
              muxOutConnector[50] = fifoOut[16][4];
              muxOutConnector[51] = fifoOut[17][4];
       end
       2: begin
              muxOutConnector[0] = fifoOut[29][7];
              muxOutConnector[1] = fifoOut[30][7];
              muxOutConnector[2] = fifoOut[31][7];
              muxOutConnector[3] = fifoOut[32][7];
              muxOutConnector[4] = fifoOut[33][7];
              muxOutConnector[5] = fifoOut[34][7];
              muxOutConnector[6] = fifoOut[35][7];
              muxOutConnector[7] = fifoOut[36][7];
              muxOutConnector[8] = fifoOut[37][7];
              muxOutConnector[9] = fifoOut[38][7];
              muxOutConnector[10] = fifoOut[39][7];
              muxOutConnector[11] = fifoOut[40][7];
              muxOutConnector[12] = fifoOut[41][7];
              muxOutConnector[13] = fifoOut[42][7];
              muxOutConnector[14] = fifoOut[43][7];
              muxOutConnector[15] = fifoOut[44][7];
              muxOutConnector[16] = fifoOut[45][7];
              muxOutConnector[17] = fifoOut[46][7];
              muxOutConnector[18] = fifoOut[47][7];
              muxOutConnector[19] = fifoOut[48][7];
              muxOutConnector[20] = fifoOut[49][7];
              muxOutConnector[21] = fifoOut[50][7];
              muxOutConnector[22] = fifoOut[51][7];
              muxOutConnector[23] = fifoOut[26][6];
              muxOutConnector[24] = fifoOut[27][6];
              muxOutConnector[25] = fifoOut[28][6];
              muxOutConnector[26] = fifoOut[18][5];
              muxOutConnector[27] = fifoOut[19][5];
              muxOutConnector[28] = fifoOut[20][5];
              muxOutConnector[29] = fifoOut[21][5];
              muxOutConnector[30] = fifoOut[22][5];
              muxOutConnector[31] = fifoOut[23][5];
              muxOutConnector[32] = fifoOut[24][5];
              muxOutConnector[33] = fifoOut[25][5];
              muxOutConnector[34] = fifoOut[0][4];
              muxOutConnector[35] = fifoOut[1][4];
              muxOutConnector[36] = fifoOut[2][4];
              muxOutConnector[37] = fifoOut[3][4];
              muxOutConnector[38] = fifoOut[4][4];
              muxOutConnector[39] = fifoOut[5][4];
              muxOutConnector[40] = fifoOut[6][4];
              muxOutConnector[41] = fifoOut[7][4];
              muxOutConnector[42] = fifoOut[8][4];
              muxOutConnector[43] = fifoOut[9][4];
              muxOutConnector[44] = fifoOut[10][4];
              muxOutConnector[45] = fifoOut[11][4];
              muxOutConnector[46] = fifoOut[12][4];
              muxOutConnector[47] = fifoOut[13][4];
              muxOutConnector[48] = fifoOut[14][4];
              muxOutConnector[49] = fifoOut[15][4];
              muxOutConnector[50] = fifoOut[16][4];
              muxOutConnector[51] = fifoOut[17][4];
       end
       3: begin
              muxOutConnector[0] = fifoOut[29][7];
              muxOutConnector[1] = fifoOut[30][7];
              muxOutConnector[2] = fifoOut[31][7];
              muxOutConnector[3] = fifoOut[32][7];
              muxOutConnector[4] = fifoOut[33][7];
              muxOutConnector[5] = fifoOut[34][7];
              muxOutConnector[6] = fifoOut[35][7];
              muxOutConnector[7] = fifoOut[36][7];
              muxOutConnector[8] = fifoOut[37][7];
              muxOutConnector[9] = fifoOut[38][7];
              muxOutConnector[10] = fifoOut[39][7];
              muxOutConnector[11] = fifoOut[40][7];
              muxOutConnector[12] = fifoOut[41][7];
              muxOutConnector[13] = fifoOut[42][7];
              muxOutConnector[14] = fifoOut[43][7];
              muxOutConnector[15] = fifoOut[44][7];
              muxOutConnector[16] = fifoOut[45][7];
              muxOutConnector[17] = fifoOut[46][7];
              muxOutConnector[18] = fifoOut[47][7];
              muxOutConnector[19] = fifoOut[48][7];
              muxOutConnector[20] = fifoOut[49][7];
              muxOutConnector[21] = fifoOut[50][7];
              muxOutConnector[22] = fifoOut[51][7];
              muxOutConnector[23] = fifoOut[26][6];
              muxOutConnector[24] = fifoOut[27][6];
              muxOutConnector[25] = fifoOut[28][6];
              muxOutConnector[26] = fifoOut[18][5];
              muxOutConnector[27] = fifoOut[19][5];
              muxOutConnector[28] = fifoOut[20][5];
              muxOutConnector[29] = fifoOut[21][5];
              muxOutConnector[30] = fifoOut[22][5];
              muxOutConnector[31] = fifoOut[23][5];
              muxOutConnector[32] = fifoOut[24][5];
              muxOutConnector[33] = fifoOut[25][5];
              muxOutConnector[34] = fifoOut[0][4];
              muxOutConnector[35] = fifoOut[1][4];
              muxOutConnector[36] = fifoOut[2][4];
              muxOutConnector[37] = fifoOut[3][4];
              muxOutConnector[38] = fifoOut[4][4];
              muxOutConnector[39] = fifoOut[5][4];
              muxOutConnector[40] = fifoOut[6][4];
              muxOutConnector[41] = fifoOut[7][4];
              muxOutConnector[42] = fifoOut[8][4];
              muxOutConnector[43] = fifoOut[9][4];
              muxOutConnector[44] = fifoOut[10][4];
              muxOutConnector[45] = fifoOut[11][4];
              muxOutConnector[46] = fifoOut[12][4];
              muxOutConnector[47] = fifoOut[13][4];
              muxOutConnector[48] = fifoOut[14][4];
              muxOutConnector[49] = fifoOut[15][4];
              muxOutConnector[50] = fifoOut[16][4];
              muxOutConnector[51] = fifoOut[17][4];
       end
       4: begin
              muxOutConnector[0] = fifoOut[29][7];
              muxOutConnector[1] = fifoOut[30][7];
              muxOutConnector[2] = fifoOut[31][7];
              muxOutConnector[3] = fifoOut[32][7];
              muxOutConnector[4] = fifoOut[33][7];
              muxOutConnector[5] = fifoOut[34][7];
              muxOutConnector[6] = fifoOut[35][7];
              muxOutConnector[7] = fifoOut[36][7];
              muxOutConnector[8] = fifoOut[37][7];
              muxOutConnector[9] = fifoOut[38][7];
              muxOutConnector[10] = fifoOut[39][7];
              muxOutConnector[11] = fifoOut[40][7];
              muxOutConnector[12] = fifoOut[41][7];
              muxOutConnector[13] = fifoOut[42][7];
              muxOutConnector[14] = fifoOut[43][7];
              muxOutConnector[15] = fifoOut[44][7];
              muxOutConnector[16] = fifoOut[45][7];
              muxOutConnector[17] = fifoOut[46][7];
              muxOutConnector[18] = fifoOut[47][7];
              muxOutConnector[19] = fifoOut[48][7];
              muxOutConnector[20] = fifoOut[49][7];
              muxOutConnector[21] = fifoOut[50][7];
              muxOutConnector[22] = fifoOut[51][7];
              muxOutConnector[23] = fifoOut[26][6];
              muxOutConnector[24] = fifoOut[27][6];
              muxOutConnector[25] = fifoOut[28][6];
              muxOutConnector[26] = fifoOut[18][5];
              muxOutConnector[27] = fifoOut[19][5];
              muxOutConnector[28] = fifoOut[20][5];
              muxOutConnector[29] = fifoOut[21][5];
              muxOutConnector[30] = fifoOut[22][5];
              muxOutConnector[31] = fifoOut[23][5];
              muxOutConnector[32] = fifoOut[24][5];
              muxOutConnector[33] = fifoOut[25][5];
              muxOutConnector[34] = fifoOut[0][4];
              muxOutConnector[35] = fifoOut[1][4];
              muxOutConnector[36] = fifoOut[2][4];
              muxOutConnector[37] = fifoOut[3][4];
              muxOutConnector[38] = fifoOut[4][4];
              muxOutConnector[39] = fifoOut[5][4];
              muxOutConnector[40] = fifoOut[6][4];
              muxOutConnector[41] = fifoOut[7][4];
              muxOutConnector[42] = fifoOut[8][4];
              muxOutConnector[43] = fifoOut[9][4];
              muxOutConnector[44] = fifoOut[10][4];
              muxOutConnector[45] = fifoOut[11][4];
              muxOutConnector[46] = fifoOut[12][4];
              muxOutConnector[47] = fifoOut[13][4];
              muxOutConnector[48] = fifoOut[14][4];
              muxOutConnector[49] = fifoOut[15][4];
              muxOutConnector[50] = fifoOut[16][4];
              muxOutConnector[51] = fifoOut[30][2];
       end
       5: begin
              muxOutConnector[0] = fifoOut[29][7];
              muxOutConnector[1] = fifoOut[30][7];
              muxOutConnector[2] = fifoOut[31][7];
              muxOutConnector[3] = fifoOut[32][7];
              muxOutConnector[4] = fifoOut[33][7];
              muxOutConnector[5] = fifoOut[34][7];
              muxOutConnector[6] = fifoOut[35][7];
              muxOutConnector[7] = fifoOut[36][7];
              muxOutConnector[8] = fifoOut[37][7];
              muxOutConnector[9] = fifoOut[38][7];
              muxOutConnector[10] = fifoOut[39][7];
              muxOutConnector[11] = fifoOut[40][7];
              muxOutConnector[12] = fifoOut[41][7];
              muxOutConnector[13] = fifoOut[42][7];
              muxOutConnector[14] = fifoOut[43][7];
              muxOutConnector[15] = fifoOut[44][7];
              muxOutConnector[16] = fifoOut[45][7];
              muxOutConnector[17] = fifoOut[46][7];
              muxOutConnector[18] = fifoOut[47][7];
              muxOutConnector[19] = fifoOut[48][7];
              muxOutConnector[20] = fifoOut[49][7];
              muxOutConnector[21] = fifoOut[50][7];
              muxOutConnector[22] = fifoOut[51][7];
              muxOutConnector[23] = fifoOut[26][6];
              muxOutConnector[24] = fifoOut[27][6];
              muxOutConnector[25] = fifoOut[28][6];
              muxOutConnector[26] = fifoOut[31][3];
              muxOutConnector[27] = fifoOut[32][3];
              muxOutConnector[28] = fifoOut[33][3];
              muxOutConnector[29] = fifoOut[34][3];
              muxOutConnector[30] = fifoOut[35][3];
              muxOutConnector[31] = fifoOut[36][3];
              muxOutConnector[32] = fifoOut[37][3];
              muxOutConnector[33] = fifoOut[38][3];
              muxOutConnector[34] = fifoOut[39][3];
              muxOutConnector[35] = fifoOut[40][3];
              muxOutConnector[36] = fifoOut[41][3];
              muxOutConnector[37] = fifoOut[42][3];
              muxOutConnector[38] = fifoOut[43][3];
              muxOutConnector[39] = fifoOut[44][3];
              muxOutConnector[40] = fifoOut[45][3];
              muxOutConnector[41] = fifoOut[46][3];
              muxOutConnector[42] = fifoOut[47][3];
              muxOutConnector[43] = fifoOut[48][3];
              muxOutConnector[44] = fifoOut[49][3];
              muxOutConnector[45] = fifoOut[50][3];
              muxOutConnector[46] = fifoOut[51][3];
              muxOutConnector[47] = fifoOut[26][2];
              muxOutConnector[48] = fifoOut[27][2];
              muxOutConnector[49] = fifoOut[28][2];
              muxOutConnector[50] = fifoOut[29][2];
              muxOutConnector[51] = fifoOut[30][2];
       end
       6: begin
              muxOutConnector[0] = fifoOut[29][7];
              muxOutConnector[1] = fifoOut[30][7];
              muxOutConnector[2] = fifoOut[31][7];
              muxOutConnector[3] = fifoOut[32][7];
              muxOutConnector[4] = fifoOut[33][7];
              muxOutConnector[5] = fifoOut[34][7];
              muxOutConnector[6] = fifoOut[35][7];
              muxOutConnector[7] = fifoOut[36][7];
              muxOutConnector[8] = fifoOut[37][7];
              muxOutConnector[9] = fifoOut[38][7];
              muxOutConnector[10] = fifoOut[39][7];
              muxOutConnector[11] = fifoOut[40][7];
              muxOutConnector[12] = fifoOut[41][7];
              muxOutConnector[13] = fifoOut[42][7];
              muxOutConnector[14] = fifoOut[43][7];
              muxOutConnector[15] = fifoOut[44][7];
              muxOutConnector[16] = fifoOut[45][7];
              muxOutConnector[17] = fifoOut[46][7];
              muxOutConnector[18] = fifoOut[47][7];
              muxOutConnector[19] = fifoOut[48][7];
              muxOutConnector[20] = fifoOut[49][7];
              muxOutConnector[21] = fifoOut[50][7];
              muxOutConnector[22] = fifoOut[51][7];
              muxOutConnector[23] = fifoOut[26][6];
              muxOutConnector[24] = fifoOut[27][6];
              muxOutConnector[25] = fifoOut[28][6];
              muxOutConnector[26] = fifoOut[31][3];
              muxOutConnector[27] = fifoOut[32][3];
              muxOutConnector[28] = fifoOut[33][3];
              muxOutConnector[29] = fifoOut[34][3];
              muxOutConnector[30] = fifoOut[35][3];
              muxOutConnector[31] = fifoOut[36][3];
              muxOutConnector[32] = fifoOut[37][3];
              muxOutConnector[33] = fifoOut[38][3];
              muxOutConnector[34] = fifoOut[39][3];
              muxOutConnector[35] = fifoOut[40][3];
              muxOutConnector[36] = fifoOut[41][3];
              muxOutConnector[37] = fifoOut[42][3];
              muxOutConnector[38] = fifoOut[43][3];
              muxOutConnector[39] = fifoOut[44][3];
              muxOutConnector[40] = fifoOut[45][3];
              muxOutConnector[41] = fifoOut[46][3];
              muxOutConnector[42] = fifoOut[47][3];
              muxOutConnector[43] = fifoOut[48][3];
              muxOutConnector[44] = fifoOut[49][3];
              muxOutConnector[45] = fifoOut[50][3];
              muxOutConnector[46] = fifoOut[51][3];
              muxOutConnector[47] = fifoOut[26][2];
              muxOutConnector[48] = fifoOut[27][2];
              muxOutConnector[49] = fifoOut[28][2];
              muxOutConnector[50] = fifoOut[29][2];
              muxOutConnector[51] = fifoOut[30][2];
       end
       7: begin
              muxOutConnector[0] = fifoOut[29][7];
              muxOutConnector[1] = fifoOut[30][7];
              muxOutConnector[2] = fifoOut[31][7];
              muxOutConnector[3] = fifoOut[32][7];
              muxOutConnector[4] = fifoOut[33][7];
              muxOutConnector[5] = fifoOut[34][7];
              muxOutConnector[6] = fifoOut[35][7];
              muxOutConnector[7] = fifoOut[36][7];
              muxOutConnector[8] = fifoOut[37][7];
              muxOutConnector[9] = fifoOut[38][7];
              muxOutConnector[10] = fifoOut[39][7];
              muxOutConnector[11] = fifoOut[40][7];
              muxOutConnector[12] = fifoOut[41][7];
              muxOutConnector[13] = fifoOut[42][7];
              muxOutConnector[14] = fifoOut[13][6];
              muxOutConnector[15] = fifoOut[14][6];
              muxOutConnector[16] = fifoOut[15][6];
              muxOutConnector[17] = fifoOut[16][6];
              muxOutConnector[18] = fifoOut[17][6];
              muxOutConnector[19] = fifoOut[18][6];
              muxOutConnector[20] = fifoOut[19][6];
              muxOutConnector[21] = fifoOut[20][6];
              muxOutConnector[22] = fifoOut[21][6];
              muxOutConnector[23] = fifoOut[22][6];
              muxOutConnector[24] = fifoOut[23][6];
              muxOutConnector[25] = fifoOut[24][6];
              muxOutConnector[26] = fifoOut[31][3];
              muxOutConnector[27] = fifoOut[32][3];
              muxOutConnector[28] = fifoOut[33][3];
              muxOutConnector[29] = fifoOut[34][3];
              muxOutConnector[30] = fifoOut[35][3];
              muxOutConnector[31] = fifoOut[36][3];
              muxOutConnector[32] = fifoOut[37][3];
              muxOutConnector[33] = fifoOut[38][3];
              muxOutConnector[34] = fifoOut[39][3];
              muxOutConnector[35] = fifoOut[40][3];
              muxOutConnector[36] = fifoOut[41][3];
              muxOutConnector[37] = fifoOut[42][3];
              muxOutConnector[38] = fifoOut[43][3];
              muxOutConnector[39] = fifoOut[44][3];
              muxOutConnector[40] = fifoOut[45][3];
              muxOutConnector[41] = fifoOut[46][3];
              muxOutConnector[42] = fifoOut[47][3];
              muxOutConnector[43] = fifoOut[48][3];
              muxOutConnector[44] = fifoOut[49][3];
              muxOutConnector[45] = fifoOut[50][3];
              muxOutConnector[46] = fifoOut[51][3];
              muxOutConnector[47] = fifoOut[26][2];
              muxOutConnector[48] = fifoOut[27][2];
              muxOutConnector[49] = fifoOut[28][2];
              muxOutConnector[50] = fifoOut[29][2];
              muxOutConnector[51] = fifoOut[30][2];
       end
       8: begin
              muxOutConnector[0] = fifoOut[25][7];
              muxOutConnector[1] = fifoOut[0][6];
              muxOutConnector[2] = fifoOut[1][6];
              muxOutConnector[3] = fifoOut[2][6];
              muxOutConnector[4] = fifoOut[3][6];
              muxOutConnector[5] = fifoOut[4][6];
              muxOutConnector[6] = fifoOut[5][6];
              muxOutConnector[7] = fifoOut[6][6];
              muxOutConnector[8] = fifoOut[7][6];
              muxOutConnector[9] = fifoOut[8][6];
              muxOutConnector[10] = fifoOut[9][6];
              muxOutConnector[11] = fifoOut[10][6];
              muxOutConnector[12] = fifoOut[11][6];
              muxOutConnector[13] = fifoOut[12][6];
              muxOutConnector[14] = fifoOut[13][6];
              muxOutConnector[15] = fifoOut[14][6];
              muxOutConnector[16] = fifoOut[15][6];
              muxOutConnector[17] = fifoOut[16][6];
              muxOutConnector[18] = fifoOut[17][6];
              muxOutConnector[19] = fifoOut[18][6];
              muxOutConnector[20] = fifoOut[19][6];
              muxOutConnector[21] = fifoOut[20][6];
              muxOutConnector[22] = fifoOut[21][6];
              muxOutConnector[23] = fifoOut[22][6];
              muxOutConnector[24] = fifoOut[23][6];
              muxOutConnector[25] = fifoOut[24][6];
              muxOutConnector[26] = fifoOut[31][3];
              muxOutConnector[27] = fifoOut[32][3];
              muxOutConnector[28] = fifoOut[33][3];
              muxOutConnector[29] = fifoOut[34][3];
              muxOutConnector[30] = fifoOut[35][3];
              muxOutConnector[31] = fifoOut[36][3];
              muxOutConnector[32] = fifoOut[37][3];
              muxOutConnector[33] = fifoOut[38][3];
              muxOutConnector[34] = fifoOut[39][3];
              muxOutConnector[35] = fifoOut[40][3];
              muxOutConnector[36] = fifoOut[41][3];
              muxOutConnector[37] = fifoOut[42][3];
              muxOutConnector[38] = fifoOut[43][3];
              muxOutConnector[39] = fifoOut[44][3];
              muxOutConnector[40] = fifoOut[45][3];
              muxOutConnector[41] = fifoOut[46][3];
              muxOutConnector[42] = fifoOut[47][3];
              muxOutConnector[43] = fifoOut[48][3];
              muxOutConnector[44] = fifoOut[49][3];
              muxOutConnector[45] = fifoOut[50][3];
              muxOutConnector[46] = fifoOut[51][3];
              muxOutConnector[47] = fifoOut[26][2];
              muxOutConnector[48] = fifoOut[27][2];
              muxOutConnector[49] = fifoOut[28][2];
              muxOutConnector[50] = fifoOut[29][2];
              muxOutConnector[51] = fifoOut[30][2];
       end
       9: begin
              muxOutConnector[0] = fifoOut[25][7];
              muxOutConnector[1] = fifoOut[0][6];
              muxOutConnector[2] = fifoOut[1][6];
              muxOutConnector[3] = fifoOut[2][6];
              muxOutConnector[4] = fifoOut[3][6];
              muxOutConnector[5] = fifoOut[4][6];
              muxOutConnector[6] = fifoOut[5][6];
              muxOutConnector[7] = fifoOut[6][6];
              muxOutConnector[8] = fifoOut[7][6];
              muxOutConnector[9] = fifoOut[8][6];
              muxOutConnector[10] = fifoOut[9][6];
              muxOutConnector[11] = fifoOut[10][6];
              muxOutConnector[12] = fifoOut[11][6];
              muxOutConnector[13] = fifoOut[12][6];
              muxOutConnector[14] = fifoOut[13][6];
              muxOutConnector[15] = fifoOut[14][6];
              muxOutConnector[16] = fifoOut[15][6];
              muxOutConnector[17] = fifoOut[16][6];
              muxOutConnector[18] = fifoOut[17][6];
              muxOutConnector[19] = fifoOut[18][6];
              muxOutConnector[20] = fifoOut[19][6];
              muxOutConnector[21] = fifoOut[20][6];
              muxOutConnector[22] = fifoOut[21][6];
              muxOutConnector[23] = fifoOut[22][6];
              muxOutConnector[24] = fifoOut[23][6];
              muxOutConnector[25] = fifoOut[24][6];
              muxOutConnector[26] = fifoOut[31][3];
              muxOutConnector[27] = fifoOut[32][3];
              muxOutConnector[28] = fifoOut[33][3];
              muxOutConnector[29] = fifoOut[34][3];
              muxOutConnector[30] = fifoOut[35][3];
              muxOutConnector[31] = fifoOut[36][3];
              muxOutConnector[32] = fifoOut[37][3];
              muxOutConnector[33] = fifoOut[38][3];
              muxOutConnector[34] = fifoOut[39][3];
              muxOutConnector[35] = fifoOut[40][3];
              muxOutConnector[36] = fifoOut[41][3];
              muxOutConnector[37] = fifoOut[42][3];
              muxOutConnector[38] = fifoOut[43][3];
              muxOutConnector[39] = fifoOut[44][3];
              muxOutConnector[40] = fifoOut[45][3];
              muxOutConnector[41] = fifoOut[46][3];
              muxOutConnector[42] = fifoOut[47][3];
              muxOutConnector[43] = fifoOut[48][3];
              muxOutConnector[44] = fifoOut[49][3];
              muxOutConnector[45] = fifoOut[50][3];
              muxOutConnector[46] = fifoOut[51][3];
              muxOutConnector[47] = fifoOut[26][2];
              muxOutConnector[48] = fifoOut[27][2];
              muxOutConnector[49] = fifoOut[28][2];
              muxOutConnector[50] = fifoOut[29][2];
              muxOutConnector[51] = fifoOut[30][2];
       end
       10: begin
              muxOutConnector[0] = fifoOut[25][7];
              muxOutConnector[1] = fifoOut[0][6];
              muxOutConnector[2] = fifoOut[1][6];
              muxOutConnector[3] = fifoOut[2][6];
              muxOutConnector[4] = fifoOut[3][6];
              muxOutConnector[5] = fifoOut[4][6];
              muxOutConnector[6] = fifoOut[5][6];
              muxOutConnector[7] = fifoOut[6][6];
              muxOutConnector[8] = fifoOut[7][6];
              muxOutConnector[9] = fifoOut[8][6];
              muxOutConnector[10] = fifoOut[9][6];
              muxOutConnector[11] = fifoOut[10][6];
              muxOutConnector[12] = fifoOut[11][6];
              muxOutConnector[13] = fifoOut[12][6];
              muxOutConnector[14] = fifoOut[13][6];
              muxOutConnector[15] = fifoOut[14][6];
              muxOutConnector[16] = fifoOut[15][6];
              muxOutConnector[17] = fifoOut[16][6];
              muxOutConnector[18] = fifoOut[17][6];
              muxOutConnector[19] = fifoOut[18][6];
              muxOutConnector[20] = fifoOut[19][6];
              muxOutConnector[21] = fifoOut[20][6];
              muxOutConnector[22] = fifoOut[21][6];
              muxOutConnector[23] = fifoOut[22][6];
              muxOutConnector[24] = fifoOut[23][6];
              muxOutConnector[25] = fifoOut[24][6];
              muxOutConnector[26] = fifoOut[31][3];
              muxOutConnector[27] = fifoOut[32][3];
              muxOutConnector[28] = fifoOut[33][3];
              muxOutConnector[29] = fifoOut[34][3];
              muxOutConnector[30] = fifoOut[35][3];
              muxOutConnector[31] = fifoOut[36][3];
              muxOutConnector[32] = fifoOut[37][3];
              muxOutConnector[33] = fifoOut[38][3];
              muxOutConnector[34] = fifoOut[39][3];
              muxOutConnector[35] = fifoOut[40][3];
              muxOutConnector[36] = fifoOut[41][3];
              muxOutConnector[37] = fifoOut[42][3];
              muxOutConnector[38] = fifoOut[43][3];
              muxOutConnector[39] = fifoOut[44][3];
              muxOutConnector[40] = fifoOut[45][3];
              muxOutConnector[41] = fifoOut[46][3];
              muxOutConnector[42] = fifoOut[47][3];
              muxOutConnector[43] = fifoOut[48][3];
              muxOutConnector[44] = fifoOut[49][3];
              muxOutConnector[45] = fifoOut[50][3];
              muxOutConnector[46] = fifoOut[51][3];
              muxOutConnector[47] = fifoOut[26][2];
              muxOutConnector[48] = fifoOut[27][2];
              muxOutConnector[49] = fifoOut[28][2];
              muxOutConnector[50] = fifoOut[29][2];
              muxOutConnector[51] = fifoOut[30][2];
       end
       11: begin
              muxOutConnector[0] = fifoOut[25][7];
              muxOutConnector[1] = fifoOut[0][6];
              muxOutConnector[2] = fifoOut[1][6];
              muxOutConnector[3] = fifoOut[2][6];
              muxOutConnector[4] = fifoOut[3][6];
              muxOutConnector[5] = fifoOut[4][6];
              muxOutConnector[6] = fifoOut[5][6];
              muxOutConnector[7] = fifoOut[6][6];
              muxOutConnector[8] = fifoOut[7][6];
              muxOutConnector[9] = fifoOut[8][6];
              muxOutConnector[10] = fifoOut[9][6];
              muxOutConnector[11] = fifoOut[10][6];
              muxOutConnector[12] = fifoOut[11][6];
              muxOutConnector[13] = fifoOut[12][6];
              muxOutConnector[14] = fifoOut[13][6];
              muxOutConnector[15] = fifoOut[14][6];
              muxOutConnector[16] = fifoOut[15][6];
              muxOutConnector[17] = fifoOut[16][6];
              muxOutConnector[18] = fifoOut[17][6];
              muxOutConnector[19] = fifoOut[18][6];
              muxOutConnector[20] = fifoOut[19][6];
              muxOutConnector[21] = fifoOut[20][6];
              muxOutConnector[22] = fifoOut[21][6];
              muxOutConnector[23] = fifoOut[22][6];
              muxOutConnector[24] = fifoOut[23][6];
              muxOutConnector[25] = fifoOut[24][6];
              muxOutConnector[26] = fifoOut[31][3];
              muxOutConnector[27] = fifoOut[32][3];
              muxOutConnector[28] = fifoOut[33][3];
              muxOutConnector[29] = fifoOut[34][3];
              muxOutConnector[30] = fifoOut[35][3];
              muxOutConnector[31] = fifoOut[36][3];
              muxOutConnector[32] = fifoOut[37][3];
              muxOutConnector[33] = fifoOut[38][3];
              muxOutConnector[34] = fifoOut[39][3];
              muxOutConnector[35] = fifoOut[40][3];
              muxOutConnector[36] = fifoOut[41][3];
              muxOutConnector[37] = fifoOut[42][3];
              muxOutConnector[38] = fifoOut[43][3];
              muxOutConnector[39] = fifoOut[44][3];
              muxOutConnector[40] = fifoOut[45][3];
              muxOutConnector[41] = fifoOut[46][3];
              muxOutConnector[42] = fifoOut[47][3];
              muxOutConnector[43] = fifoOut[48][3];
              muxOutConnector[44] = fifoOut[49][3];
              muxOutConnector[45] = fifoOut[50][3];
              muxOutConnector[46] = fifoOut[51][3];
              muxOutConnector[47] = fifoOut[26][2];
              muxOutConnector[48] = fifoOut[27][2];
              muxOutConnector[49] = fifoOut[28][2];
              muxOutConnector[50] = fifoOut[29][2];
              muxOutConnector[51] = fifoOut[30][2];
       end
       12: begin
              muxOutConnector[0] = fifoOut[25][7];
              muxOutConnector[1] = fifoOut[0][6];
              muxOutConnector[2] = fifoOut[1][6];
              muxOutConnector[3] = fifoOut[2][6];
              muxOutConnector[4] = fifoOut[3][6];
              muxOutConnector[5] = fifoOut[4][6];
              muxOutConnector[6] = fifoOut[5][6];
              muxOutConnector[7] = fifoOut[6][6];
              muxOutConnector[8] = fifoOut[7][6];
              muxOutConnector[9] = fifoOut[8][6];
              muxOutConnector[10] = fifoOut[9][6];
              muxOutConnector[11] = fifoOut[10][6];
              muxOutConnector[12] = fifoOut[11][6];
              muxOutConnector[13] = fifoOut[12][6];
              muxOutConnector[14] = fifoOut[13][6];
              muxOutConnector[15] = fifoOut[14][6];
              muxOutConnector[16] = fifoOut[15][6];
              muxOutConnector[17] = fifoOut[16][6];
              muxOutConnector[18] = fifoOut[17][6];
              muxOutConnector[19] = fifoOut[18][6];
              muxOutConnector[20] = fifoOut[19][6];
              muxOutConnector[21] = fifoOut[20][6];
              muxOutConnector[22] = fifoOut[21][6];
              muxOutConnector[23] = fifoOut[22][6];
              muxOutConnector[24] = fifoOut[23][6];
              muxOutConnector[25] = fifoOut[24][6];
              muxOutConnector[26] = fifoOut[31][3];
              muxOutConnector[27] = fifoOut[32][3];
              muxOutConnector[28] = fifoOut[33][3];
              muxOutConnector[29] = fifoOut[34][3];
              muxOutConnector[30] = fifoOut[35][3];
              muxOutConnector[31] = fifoOut[36][3];
              muxOutConnector[32] = fifoOut[37][3];
              muxOutConnector[33] = fifoOut[38][3];
              muxOutConnector[34] = fifoOut[39][3];
              muxOutConnector[35] = fifoOut[40][3];
              muxOutConnector[36] = fifoOut[41][3];
              muxOutConnector[37] = fifoOut[42][3];
              muxOutConnector[38] = fifoOut[43][3];
              muxOutConnector[39] = fifoOut[44][3];
              muxOutConnector[40] = fifoOut[45][3];
              muxOutConnector[41] = fifoOut[46][3];
              muxOutConnector[42] = fifoOut[47][3];
              muxOutConnector[43] = fifoOut[48][3];
              muxOutConnector[44] = fifoOut[49][3];
              muxOutConnector[45] = fifoOut[50][3];
              muxOutConnector[46] = fifoOut[51][3];
              muxOutConnector[47] = fifoOut[26][2];
              muxOutConnector[48] = fifoOut[27][2];
              muxOutConnector[49] = fifoOut[28][2];
              muxOutConnector[50] = fifoOut[29][2];
              muxOutConnector[51] = fifoOut[30][2];
       end
       13: begin
              muxOutConnector[0] = fifoOut[25][7];
              muxOutConnector[1] = fifoOut[0][6];
              muxOutConnector[2] = fifoOut[1][6];
              muxOutConnector[3] = fifoOut[2][6];
              muxOutConnector[4] = fifoOut[3][6];
              muxOutConnector[5] = fifoOut[4][6];
              muxOutConnector[6] = fifoOut[5][6];
              muxOutConnector[7] = fifoOut[6][6];
              muxOutConnector[8] = fifoOut[7][6];
              muxOutConnector[9] = fifoOut[8][6];
              muxOutConnector[10] = fifoOut[9][6];
              muxOutConnector[11] = fifoOut[10][6];
              muxOutConnector[12] = fifoOut[11][6];
              muxOutConnector[13] = fifoOut[12][6];
              muxOutConnector[14] = fifoOut[13][6];
              muxOutConnector[15] = fifoOut[14][6];
              muxOutConnector[16] = fifoOut[15][6];
              muxOutConnector[17] = fifoOut[16][6];
              muxOutConnector[18] = fifoOut[17][6];
              muxOutConnector[19] = fifoOut[18][6];
              muxOutConnector[20] = fifoOut[19][6];
              muxOutConnector[21] = fifoOut[20][6];
              muxOutConnector[22] = fifoOut[21][6];
              muxOutConnector[23] = fifoOut[22][6];
              muxOutConnector[24] = fifoOut[23][6];
              muxOutConnector[25] = fifoOut[24][6];
              muxOutConnector[26] = fifoOut[31][3];
              muxOutConnector[27] = fifoOut[32][3];
              muxOutConnector[28] = fifoOut[33][3];
              muxOutConnector[29] = fifoOut[34][3];
              muxOutConnector[30] = fifoOut[35][3];
              muxOutConnector[31] = fifoOut[36][3];
              muxOutConnector[32] = fifoOut[37][3];
              muxOutConnector[33] = fifoOut[38][3];
              muxOutConnector[34] = fifoOut[39][3];
              muxOutConnector[35] = fifoOut[40][3];
              muxOutConnector[36] = fifoOut[41][3];
              muxOutConnector[37] = fifoOut[42][3];
              muxOutConnector[38] = fifoOut[43][3];
              muxOutConnector[39] = fifoOut[44][3];
              muxOutConnector[40] = fifoOut[45][3];
              muxOutConnector[41] = fifoOut[46][3];
              muxOutConnector[42] = fifoOut[47][3];
              muxOutConnector[43] = fifoOut[48][3];
              muxOutConnector[44] = fifoOut[49][3];
              muxOutConnector[45] = fifoOut[50][3];
              muxOutConnector[46] = fifoOut[51][3];
              muxOutConnector[47] = fifoOut[26][2];
              muxOutConnector[48] = fifoOut[27][2];
              muxOutConnector[49] = fifoOut[28][2];
              muxOutConnector[50] = fifoOut[29][2];
              muxOutConnector[51] = fifoOut[30][2];
       end
       14: begin
              muxOutConnector[0] = fifoOut[25][7];
              muxOutConnector[1] = fifoOut[0][6];
              muxOutConnector[2] = fifoOut[1][6];
              muxOutConnector[3] = fifoOut[2][6];
              muxOutConnector[4] = fifoOut[3][6];
              muxOutConnector[5] = fifoOut[4][6];
              muxOutConnector[6] = fifoOut[5][6];
              muxOutConnector[7] = fifoOut[6][6];
              muxOutConnector[8] = fifoOut[7][6];
              muxOutConnector[9] = fifoOut[8][6];
              muxOutConnector[10] = fifoOut[9][6];
              muxOutConnector[11] = fifoOut[10][6];
              muxOutConnector[12] = fifoOut[11][6];
              muxOutConnector[13] = fifoOut[12][6];
              muxOutConnector[14] = fifoOut[13][6];
              muxOutConnector[15] = fifoOut[14][6];
              muxOutConnector[16] = fifoOut[15][6];
              muxOutConnector[17] = fifoOut[16][6];
              muxOutConnector[18] = fifoOut[17][6];
              muxOutConnector[19] = fifoOut[18][6];
              muxOutConnector[20] = fifoOut[19][6];
              muxOutConnector[21] = fifoOut[20][6];
              muxOutConnector[22] = fifoOut[21][6];
              muxOutConnector[23] = fifoOut[22][6];
              muxOutConnector[24] = fifoOut[23][6];
              muxOutConnector[25] = fifoOut[24][6];
              muxOutConnector[26] = fifoOut[31][3];
              muxOutConnector[27] = fifoOut[32][3];
              muxOutConnector[28] = fifoOut[33][3];
              muxOutConnector[29] = fifoOut[34][3];
              muxOutConnector[30] = fifoOut[35][3];
              muxOutConnector[31] = fifoOut[36][3];
              muxOutConnector[32] = fifoOut[37][3];
              muxOutConnector[33] = fifoOut[38][3];
              muxOutConnector[34] = fifoOut[39][3];
              muxOutConnector[35] = fifoOut[40][3];
              muxOutConnector[36] = fifoOut[41][3];
              muxOutConnector[37] = fifoOut[42][3];
              muxOutConnector[38] = fifoOut[13][2];
              muxOutConnector[39] = fifoOut[14][2];
              muxOutConnector[40] = fifoOut[15][2];
              muxOutConnector[41] = fifoOut[16][2];
              muxOutConnector[42] = fifoOut[17][2];
              muxOutConnector[43] = fifoOut[18][2];
              muxOutConnector[44] = fifoOut[19][2];
              muxOutConnector[45] = fifoOut[20][2];
              muxOutConnector[46] = fifoOut[21][2];
              muxOutConnector[47] = fifoOut[22][2];
              muxOutConnector[48] = fifoOut[23][2];
              muxOutConnector[49] = fifoOut[24][2];
              muxOutConnector[50] = fifoOut[25][2];
              muxOutConnector[51] = fifoOut[0][1];
       end
       15: begin
              muxOutConnector[0] = fifoOut[25][7];
              muxOutConnector[1] = fifoOut[0][6];
              muxOutConnector[2] = fifoOut[1][6];
              muxOutConnector[3] = fifoOut[2][6];
              muxOutConnector[4] = fifoOut[3][6];
              muxOutConnector[5] = fifoOut[4][6];
              muxOutConnector[6] = fifoOut[5][6];
              muxOutConnector[7] = fifoOut[6][6];
              muxOutConnector[8] = fifoOut[7][6];
              muxOutConnector[9] = fifoOut[8][6];
              muxOutConnector[10] = fifoOut[9][6];
              muxOutConnector[11] = fifoOut[10][6];
              muxOutConnector[12] = fifoOut[11][6];
              muxOutConnector[13] = fifoOut[12][6];
              muxOutConnector[14] = fifoOut[13][6];
              muxOutConnector[15] = fifoOut[14][6];
              muxOutConnector[16] = fifoOut[15][6];
              muxOutConnector[17] = fifoOut[16][6];
              muxOutConnector[18] = fifoOut[17][6];
              muxOutConnector[19] = fifoOut[18][6];
              muxOutConnector[20] = fifoOut[19][6];
              muxOutConnector[21] = fifoOut[20][6];
              muxOutConnector[22] = fifoOut[21][6];
              muxOutConnector[23] = fifoOut[22][6];
              muxOutConnector[24] = fifoOut[23][6];
              muxOutConnector[25] = fifoOut[24][6];
              muxOutConnector[26] = fifoOut[1][2];
              muxOutConnector[27] = fifoOut[2][2];
              muxOutConnector[28] = fifoOut[3][2];
              muxOutConnector[29] = fifoOut[4][2];
              muxOutConnector[30] = fifoOut[5][2];
              muxOutConnector[31] = fifoOut[6][2];
              muxOutConnector[32] = fifoOut[7][2];
              muxOutConnector[33] = fifoOut[8][2];
              muxOutConnector[34] = fifoOut[9][2];
              muxOutConnector[35] = fifoOut[10][2];
              muxOutConnector[36] = fifoOut[11][2];
              muxOutConnector[37] = fifoOut[12][2];
              muxOutConnector[38] = fifoOut[13][2];
              muxOutConnector[39] = fifoOut[14][2];
              muxOutConnector[40] = fifoOut[15][2];
              muxOutConnector[41] = fifoOut[16][2];
              muxOutConnector[42] = fifoOut[17][2];
              muxOutConnector[43] = fifoOut[18][2];
              muxOutConnector[44] = fifoOut[19][2];
              muxOutConnector[45] = fifoOut[20][2];
              muxOutConnector[46] = fifoOut[21][2];
              muxOutConnector[47] = fifoOut[22][2];
              muxOutConnector[48] = fifoOut[23][2];
              muxOutConnector[49] = fifoOut[24][2];
              muxOutConnector[50] = fifoOut[25][2];
              muxOutConnector[51] = fifoOut[0][1];
       end
       16: begin
              muxOutConnector[0] = fifoOut[25][7];
              muxOutConnector[1] = fifoOut[0][6];
              muxOutConnector[2] = fifoOut[1][6];
              muxOutConnector[3] = fifoOut[2][6];
              muxOutConnector[4] = fifoOut[3][6];
              muxOutConnector[5] = fifoOut[4][6];
              muxOutConnector[6] = fifoOut[5][6];
              muxOutConnector[7] = fifoOut[6][6];
              muxOutConnector[8] = fifoOut[7][6];
              muxOutConnector[9] = fifoOut[8][6];
              muxOutConnector[10] = fifoOut[9][6];
              muxOutConnector[11] = fifoOut[10][6];
              muxOutConnector[12] = fifoOut[11][6];
              muxOutConnector[13] = fifoOut[12][6];
              muxOutConnector[14] = fifoOut[13][6];
              muxOutConnector[15] = fifoOut[14][6];
              muxOutConnector[16] = fifoOut[15][6];
              muxOutConnector[17] = fifoOut[16][6];
              muxOutConnector[18] = fifoOut[17][6];
              muxOutConnector[19] = fifoOut[18][6];
              muxOutConnector[20] = fifoOut[19][6];
              muxOutConnector[21] = fifoOut[20][6];
              muxOutConnector[22] = fifoOut[21][6];
              muxOutConnector[23] = fifoOut[22][6];
              muxOutConnector[24] = fifoOut[23][6];
              muxOutConnector[25] = fifoOut[24][6];
              muxOutConnector[26] = fifoOut[1][2];
              muxOutConnector[27] = fifoOut[2][2];
              muxOutConnector[28] = fifoOut[3][2];
              muxOutConnector[29] = fifoOut[4][2];
              muxOutConnector[30] = fifoOut[5][2];
              muxOutConnector[31] = fifoOut[6][2];
              muxOutConnector[32] = fifoOut[7][2];
              muxOutConnector[33] = fifoOut[8][2];
              muxOutConnector[34] = fifoOut[9][2];
              muxOutConnector[35] = fifoOut[10][2];
              muxOutConnector[36] = fifoOut[11][2];
              muxOutConnector[37] = fifoOut[12][2];
              muxOutConnector[38] = fifoOut[13][2];
              muxOutConnector[39] = fifoOut[14][2];
              muxOutConnector[40] = fifoOut[15][2];
              muxOutConnector[41] = fifoOut[16][2];
              muxOutConnector[42] = fifoOut[17][2];
              muxOutConnector[43] = fifoOut[18][2];
              muxOutConnector[44] = fifoOut[19][2];
              muxOutConnector[45] = fifoOut[20][2];
              muxOutConnector[46] = fifoOut[21][2];
              muxOutConnector[47] = fifoOut[22][2];
              muxOutConnector[48] = fifoOut[23][2];
              muxOutConnector[49] = fifoOut[24][2];
              muxOutConnector[50] = fifoOut[25][2];
              muxOutConnector[51] = fifoOut[0][1];
       end
       17: begin
              muxOutConnector[0] = fifoOut[25][7];
              muxOutConnector[1] = fifoOut[0][6];
              muxOutConnector[2] = fifoOut[1][6];
              muxOutConnector[3] = fifoOut[2][6];
              muxOutConnector[4] = fifoOut[3][6];
              muxOutConnector[5] = fifoOut[4][6];
              muxOutConnector[6] = fifoOut[5][6];
              muxOutConnector[7] = fifoOut[6][6];
              muxOutConnector[8] = fifoOut[7][6];
              muxOutConnector[9] = fifoOut[8][6];
              muxOutConnector[10] = fifoOut[9][6];
              muxOutConnector[11] = fifoOut[10][6];
              muxOutConnector[12] = fifoOut[11][6];
              muxOutConnector[13] = fifoOut[12][6];
              muxOutConnector[14] = fifoOut[13][6];
              muxOutConnector[15] = fifoOut[14][6];
              muxOutConnector[16] = fifoOut[15][6];
              muxOutConnector[17] = fifoOut[16][6];
              muxOutConnector[18] = fifoOut[30][4];
              muxOutConnector[19] = fifoOut[31][4];
              muxOutConnector[20] = fifoOut[32][4];
              muxOutConnector[21] = fifoOut[33][4];
              muxOutConnector[22] = fifoOut[34][4];
              muxOutConnector[23] = fifoOut[35][4];
              muxOutConnector[24] = fifoOut[36][4];
              muxOutConnector[25] = fifoOut[37][4];
              muxOutConnector[26] = fifoOut[1][2];
              muxOutConnector[27] = fifoOut[2][2];
              muxOutConnector[28] = fifoOut[3][2];
              muxOutConnector[29] = fifoOut[4][2];
              muxOutConnector[30] = fifoOut[5][2];
              muxOutConnector[31] = fifoOut[6][2];
              muxOutConnector[32] = fifoOut[7][2];
              muxOutConnector[33] = fifoOut[8][2];
              muxOutConnector[34] = fifoOut[9][2];
              muxOutConnector[35] = fifoOut[10][2];
              muxOutConnector[36] = fifoOut[11][2];
              muxOutConnector[37] = fifoOut[12][2];
              muxOutConnector[38] = fifoOut[13][2];
              muxOutConnector[39] = fifoOut[14][2];
              muxOutConnector[40] = fifoOut[15][2];
              muxOutConnector[41] = fifoOut[16][2];
              muxOutConnector[42] = fifoOut[17][2];
              muxOutConnector[43] = fifoOut[18][2];
              muxOutConnector[44] = fifoOut[19][2];
              muxOutConnector[45] = fifoOut[20][2];
              muxOutConnector[46] = fifoOut[21][2];
              muxOutConnector[47] = fifoOut[22][2];
              muxOutConnector[48] = fifoOut[23][2];
              muxOutConnector[49] = fifoOut[24][2];
              muxOutConnector[50] = fifoOut[25][2];
              muxOutConnector[51] = fifoOut[0][1];
       end
       18: begin
              muxOutConnector[0] = fifoOut[38][5];
              muxOutConnector[1] = fifoOut[39][5];
              muxOutConnector[2] = fifoOut[40][5];
              muxOutConnector[3] = fifoOut[41][5];
              muxOutConnector[4] = fifoOut[42][5];
              muxOutConnector[5] = fifoOut[43][5];
              muxOutConnector[6] = fifoOut[44][5];
              muxOutConnector[7] = fifoOut[45][5];
              muxOutConnector[8] = fifoOut[46][5];
              muxOutConnector[9] = fifoOut[47][5];
              muxOutConnector[10] = fifoOut[48][5];
              muxOutConnector[11] = fifoOut[49][5];
              muxOutConnector[12] = fifoOut[50][5];
              muxOutConnector[13] = fifoOut[51][5];
              muxOutConnector[14] = fifoOut[26][4];
              muxOutConnector[15] = fifoOut[27][4];
              muxOutConnector[16] = fifoOut[28][4];
              muxOutConnector[17] = fifoOut[29][4];
              muxOutConnector[18] = fifoOut[30][4];
              muxOutConnector[19] = fifoOut[31][4];
              muxOutConnector[20] = fifoOut[32][4];
              muxOutConnector[21] = fifoOut[33][4];
              muxOutConnector[22] = fifoOut[34][4];
              muxOutConnector[23] = fifoOut[35][4];
              muxOutConnector[24] = fifoOut[36][4];
              muxOutConnector[25] = fifoOut[37][4];
              muxOutConnector[26] = fifoOut[1][2];
              muxOutConnector[27] = fifoOut[2][2];
              muxOutConnector[28] = fifoOut[3][2];
              muxOutConnector[29] = fifoOut[4][2];
              muxOutConnector[30] = fifoOut[5][2];
              muxOutConnector[31] = fifoOut[6][2];
              muxOutConnector[32] = fifoOut[7][2];
              muxOutConnector[33] = fifoOut[8][2];
              muxOutConnector[34] = fifoOut[9][2];
              muxOutConnector[35] = fifoOut[10][2];
              muxOutConnector[36] = fifoOut[11][2];
              muxOutConnector[37] = fifoOut[12][2];
              muxOutConnector[38] = fifoOut[13][2];
              muxOutConnector[39] = fifoOut[14][2];
              muxOutConnector[40] = fifoOut[15][2];
              muxOutConnector[41] = fifoOut[16][2];
              muxOutConnector[42] = fifoOut[17][2];
              muxOutConnector[43] = fifoOut[18][2];
              muxOutConnector[44] = fifoOut[19][2];
              muxOutConnector[45] = fifoOut[20][2];
              muxOutConnector[46] = fifoOut[21][2];
              muxOutConnector[47] = fifoOut[22][2];
              muxOutConnector[48] = fifoOut[23][2];
              muxOutConnector[49] = fifoOut[24][2];
              muxOutConnector[50] = fifoOut[25][2];
              muxOutConnector[51] = fifoOut[0][1];
       end
       19: begin
              muxOutConnector[0] = fifoOut[38][5];
              muxOutConnector[1] = fifoOut[39][5];
              muxOutConnector[2] = fifoOut[40][5];
              muxOutConnector[3] = fifoOut[41][5];
              muxOutConnector[4] = fifoOut[42][5];
              muxOutConnector[5] = fifoOut[43][5];
              muxOutConnector[6] = fifoOut[44][5];
              muxOutConnector[7] = fifoOut[45][5];
              muxOutConnector[8] = fifoOut[46][5];
              muxOutConnector[9] = fifoOut[47][5];
              muxOutConnector[10] = fifoOut[48][5];
              muxOutConnector[11] = fifoOut[49][5];
              muxOutConnector[12] = fifoOut[50][5];
              muxOutConnector[13] = fifoOut[51][5];
              muxOutConnector[14] = fifoOut[26][4];
              muxOutConnector[15] = fifoOut[27][4];
              muxOutConnector[16] = fifoOut[28][4];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[1][2];
              muxOutConnector[27] = fifoOut[2][2];
              muxOutConnector[28] = fifoOut[3][2];
              muxOutConnector[29] = fifoOut[4][2];
              muxOutConnector[30] = fifoOut[5][2];
              muxOutConnector[31] = fifoOut[6][2];
              muxOutConnector[32] = fifoOut[7][2];
              muxOutConnector[33] = fifoOut[8][2];
              muxOutConnector[34] = fifoOut[9][2];
              muxOutConnector[35] = fifoOut[10][2];
              muxOutConnector[36] = fifoOut[11][2];
              muxOutConnector[37] = fifoOut[12][2];
              muxOutConnector[38] = fifoOut[13][2];
              muxOutConnector[39] = fifoOut[14][2];
              muxOutConnector[40] = fifoOut[15][2];
              muxOutConnector[41] = fifoOut[16][2];
              muxOutConnector[42] = fifoOut[17][2];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
