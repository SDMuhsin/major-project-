`timescale 1ns / 1ps
module LMem1To0_511_circ9_combined_ys_yu_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        rxIn,
        load_input_en,
        iteration_0_indicator,
        feedback_en,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter r_lower = 32;
parameter c = 17;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input load_input_en;
input iteration_0_indicator;
input [ADDRESSWIDTH-1:0]unloadAddress;
input feedback_en;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input [ r_lower * w - 1 : 0 ] rxIn; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
wire [w-1:0]rxInConnector[r_lower-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

generate
    for (k=0;k<r_lower;k=k+1)begin:assign_rx
        assign rxInConnector[k] = rxIn[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            if(feedback_en)begin
                 fifoOut[i][0] <= fifoOut[i][c-1];
            end
            else if(load_input_en)begin
                 if(i < r_lower)begin
                   fifoOut[i][0] = rxInConnector[i];
                 end
                 else begin
                   fifoOut[i][0] = maxVal;
                 end
            end
            else begin
                 fifoOut[i][0] <= ly0InConnector[i];
            end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
       0: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = fifoOut[1][11][w-1];
              unloadMuxOut[24] = fifoOut[2][11][w-1];
              unloadMuxOut[25] = fifoOut[3][11][w-1];
              unloadMuxOut[26] = fifoOut[4][11][w-1];
              unloadMuxOut[27] = fifoOut[5][11][w-1];
              unloadMuxOut[28] = fifoOut[6][11][w-1];
              unloadMuxOut[29] = fifoOut[7][11][w-1];
              unloadMuxOut[30] = fifoOut[8][11][w-1];
              unloadMuxOut[31] = fifoOut[9][11][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[10][12][w-1];
              unloadMuxOut[1] = fifoOut[11][12][w-1];
              unloadMuxOut[2] = fifoOut[12][12][w-1];
              unloadMuxOut[3] = fifoOut[13][12][w-1];
              unloadMuxOut[4] = fifoOut[14][12][w-1];
              unloadMuxOut[5] = fifoOut[15][12][w-1];
              unloadMuxOut[6] = fifoOut[16][12][w-1];
              unloadMuxOut[7] = fifoOut[17][12][w-1];
              unloadMuxOut[8] = fifoOut[18][12][w-1];
              unloadMuxOut[9] = fifoOut[19][12][w-1];
              unloadMuxOut[10] = fifoOut[20][12][w-1];
              unloadMuxOut[11] = fifoOut[21][12][w-1];
              unloadMuxOut[12] = fifoOut[22][12][w-1];
              unloadMuxOut[13] = fifoOut[23][12][w-1];
              unloadMuxOut[14] = fifoOut[24][12][w-1];
              unloadMuxOut[15] = fifoOut[25][12][w-1];
              unloadMuxOut[16] = fifoOut[0][11][w-1];
              unloadMuxOut[17] = fifoOut[1][11][w-1];
              unloadMuxOut[18] = fifoOut[2][11][w-1];
              unloadMuxOut[19] = fifoOut[3][11][w-1];
              unloadMuxOut[20] = fifoOut[4][11][w-1];
              unloadMuxOut[21] = fifoOut[5][11][w-1];
              unloadMuxOut[22] = fifoOut[6][11][w-1];
              unloadMuxOut[23] = fifoOut[7][11][w-1];
              unloadMuxOut[24] = fifoOut[8][11][w-1];
              unloadMuxOut[25] = fifoOut[9][11][w-1];
              unloadMuxOut[26] = fifoOut[10][11][w-1];
              unloadMuxOut[27] = fifoOut[11][11][w-1];
              unloadMuxOut[28] = fifoOut[12][11][w-1];
              unloadMuxOut[29] = fifoOut[13][11][w-1];
              unloadMuxOut[30] = fifoOut[14][11][w-1];
              unloadMuxOut[31] = fifoOut[15][11][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[16][12][w-1];
              unloadMuxOut[1] = fifoOut[17][12][w-1];
              unloadMuxOut[2] = fifoOut[18][12][w-1];
              unloadMuxOut[3] = fifoOut[19][12][w-1];
              unloadMuxOut[4] = fifoOut[20][12][w-1];
              unloadMuxOut[5] = fifoOut[21][12][w-1];
              unloadMuxOut[6] = fifoOut[22][12][w-1];
              unloadMuxOut[7] = fifoOut[23][12][w-1];
              unloadMuxOut[8] = fifoOut[24][12][w-1];
              unloadMuxOut[9] = fifoOut[25][12][w-1];
              unloadMuxOut[10] = fifoOut[0][11][w-1];
              unloadMuxOut[11] = fifoOut[1][11][w-1];
              unloadMuxOut[12] = fifoOut[2][11][w-1];
              unloadMuxOut[13] = fifoOut[3][11][w-1];
              unloadMuxOut[14] = fifoOut[4][11][w-1];
              unloadMuxOut[15] = fifoOut[5][11][w-1];
              unloadMuxOut[16] = fifoOut[6][11][w-1];
              unloadMuxOut[17] = fifoOut[7][11][w-1];
              unloadMuxOut[18] = fifoOut[8][11][w-1];
              unloadMuxOut[19] = fifoOut[9][11][w-1];
              unloadMuxOut[20] = fifoOut[10][11][w-1];
              unloadMuxOut[21] = fifoOut[11][11][w-1];
              unloadMuxOut[22] = fifoOut[12][11][w-1];
              unloadMuxOut[23] = fifoOut[13][11][w-1];
              unloadMuxOut[24] = fifoOut[14][11][w-1];
              unloadMuxOut[25] = fifoOut[15][11][w-1];
              unloadMuxOut[26] = fifoOut[16][11][w-1];
              unloadMuxOut[27] = fifoOut[17][11][w-1];
              unloadMuxOut[28] = fifoOut[18][11][w-1];
              unloadMuxOut[29] = fifoOut[26][16][w-1];
              unloadMuxOut[30] = fifoOut[27][16][w-1];
              unloadMuxOut[31] = fifoOut[28][16][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[22][12][w-1];
              unloadMuxOut[1] = fifoOut[23][12][w-1];
              unloadMuxOut[2] = fifoOut[24][12][w-1];
              unloadMuxOut[3] = fifoOut[25][12][w-1];
              unloadMuxOut[4] = fifoOut[0][11][w-1];
              unloadMuxOut[5] = fifoOut[1][11][w-1];
              unloadMuxOut[6] = fifoOut[2][11][w-1];
              unloadMuxOut[7] = fifoOut[3][11][w-1];
              unloadMuxOut[8] = fifoOut[4][11][w-1];
              unloadMuxOut[9] = fifoOut[5][11][w-1];
              unloadMuxOut[10] = fifoOut[6][11][w-1];
              unloadMuxOut[11] = fifoOut[7][11][w-1];
              unloadMuxOut[12] = fifoOut[8][11][w-1];
              unloadMuxOut[13] = fifoOut[9][11][w-1];
              unloadMuxOut[14] = fifoOut[10][11][w-1];
              unloadMuxOut[15] = fifoOut[11][11][w-1];
              unloadMuxOut[16] = fifoOut[12][11][w-1];
              unloadMuxOut[17] = fifoOut[13][11][w-1];
              unloadMuxOut[18] = fifoOut[14][11][w-1];
              unloadMuxOut[19] = fifoOut[15][11][w-1];
              unloadMuxOut[20] = fifoOut[16][11][w-1];
              unloadMuxOut[21] = fifoOut[17][11][w-1];
              unloadMuxOut[22] = fifoOut[18][11][w-1];
              unloadMuxOut[23] = fifoOut[26][16][w-1];
              unloadMuxOut[24] = fifoOut[27][16][w-1];
              unloadMuxOut[25] = fifoOut[28][16][w-1];
              unloadMuxOut[26] = fifoOut[29][16][w-1];
              unloadMuxOut[27] = fifoOut[30][16][w-1];
              unloadMuxOut[28] = fifoOut[31][16][w-1];
              unloadMuxOut[29] = fifoOut[32][16][w-1];
              unloadMuxOut[30] = fifoOut[33][16][w-1];
              unloadMuxOut[31] = fifoOut[34][16][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[2][11][w-1];
              unloadMuxOut[1] = fifoOut[3][11][w-1];
              unloadMuxOut[2] = fifoOut[4][11][w-1];
              unloadMuxOut[3] = fifoOut[5][11][w-1];
              unloadMuxOut[4] = fifoOut[6][11][w-1];
              unloadMuxOut[5] = fifoOut[7][11][w-1];
              unloadMuxOut[6] = fifoOut[8][11][w-1];
              unloadMuxOut[7] = fifoOut[9][11][w-1];
              unloadMuxOut[8] = fifoOut[10][11][w-1];
              unloadMuxOut[9] = fifoOut[11][11][w-1];
              unloadMuxOut[10] = fifoOut[12][11][w-1];
              unloadMuxOut[11] = fifoOut[13][11][w-1];
              unloadMuxOut[12] = fifoOut[14][11][w-1];
              unloadMuxOut[13] = fifoOut[15][11][w-1];
              unloadMuxOut[14] = fifoOut[16][11][w-1];
              unloadMuxOut[15] = fifoOut[17][11][w-1];
              unloadMuxOut[16] = fifoOut[18][11][w-1];
              unloadMuxOut[17] = fifoOut[26][16][w-1];
              unloadMuxOut[18] = fifoOut[27][16][w-1];
              unloadMuxOut[19] = fifoOut[28][16][w-1];
              unloadMuxOut[20] = fifoOut[29][16][w-1];
              unloadMuxOut[21] = fifoOut[30][16][w-1];
              unloadMuxOut[22] = fifoOut[31][16][w-1];
              unloadMuxOut[23] = fifoOut[32][16][w-1];
              unloadMuxOut[24] = fifoOut[33][16][w-1];
              unloadMuxOut[25] = fifoOut[34][16][w-1];
              unloadMuxOut[26] = fifoOut[35][16][w-1];
              unloadMuxOut[27] = fifoOut[36][16][w-1];
              unloadMuxOut[28] = fifoOut[37][16][w-1];
              unloadMuxOut[29] = fifoOut[38][16][w-1];
              unloadMuxOut[30] = fifoOut[39][16][w-1];
              unloadMuxOut[31] = fifoOut[40][16][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[8][11][w-1];
              unloadMuxOut[1] = fifoOut[9][11][w-1];
              unloadMuxOut[2] = fifoOut[10][11][w-1];
              unloadMuxOut[3] = fifoOut[11][11][w-1];
              unloadMuxOut[4] = fifoOut[12][11][w-1];
              unloadMuxOut[5] = fifoOut[13][11][w-1];
              unloadMuxOut[6] = fifoOut[14][11][w-1];
              unloadMuxOut[7] = fifoOut[15][11][w-1];
              unloadMuxOut[8] = fifoOut[16][11][w-1];
              unloadMuxOut[9] = fifoOut[17][11][w-1];
              unloadMuxOut[10] = fifoOut[18][11][w-1];
              unloadMuxOut[11] = fifoOut[26][16][w-1];
              unloadMuxOut[12] = fifoOut[27][16][w-1];
              unloadMuxOut[13] = fifoOut[28][16][w-1];
              unloadMuxOut[14] = fifoOut[29][16][w-1];
              unloadMuxOut[15] = fifoOut[30][16][w-1];
              unloadMuxOut[16] = fifoOut[31][16][w-1];
              unloadMuxOut[17] = fifoOut[32][16][w-1];
              unloadMuxOut[18] = fifoOut[33][16][w-1];
              unloadMuxOut[19] = fifoOut[34][16][w-1];
              unloadMuxOut[20] = fifoOut[35][16][w-1];
              unloadMuxOut[21] = fifoOut[36][16][w-1];
              unloadMuxOut[22] = fifoOut[37][16][w-1];
              unloadMuxOut[23] = fifoOut[38][16][w-1];
              unloadMuxOut[24] = fifoOut[39][16][w-1];
              unloadMuxOut[25] = fifoOut[40][16][w-1];
              unloadMuxOut[26] = fifoOut[41][16][w-1];
              unloadMuxOut[27] = fifoOut[42][16][w-1];
              unloadMuxOut[28] = fifoOut[43][16][w-1];
              unloadMuxOut[29] = fifoOut[44][16][w-1];
              unloadMuxOut[30] = fifoOut[45][16][w-1];
              unloadMuxOut[31] = fifoOut[46][16][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[14][11][w-1];
              unloadMuxOut[1] = fifoOut[15][11][w-1];
              unloadMuxOut[2] = fifoOut[16][11][w-1];
              unloadMuxOut[3] = fifoOut[17][11][w-1];
              unloadMuxOut[4] = fifoOut[18][11][w-1];
              unloadMuxOut[5] = fifoOut[26][16][w-1];
              unloadMuxOut[6] = fifoOut[27][16][w-1];
              unloadMuxOut[7] = fifoOut[28][16][w-1];
              unloadMuxOut[8] = fifoOut[29][16][w-1];
              unloadMuxOut[9] = fifoOut[30][16][w-1];
              unloadMuxOut[10] = fifoOut[31][16][w-1];
              unloadMuxOut[11] = fifoOut[32][16][w-1];
              unloadMuxOut[12] = fifoOut[33][16][w-1];
              unloadMuxOut[13] = fifoOut[34][16][w-1];
              unloadMuxOut[14] = fifoOut[35][16][w-1];
              unloadMuxOut[15] = fifoOut[36][16][w-1];
              unloadMuxOut[16] = fifoOut[37][16][w-1];
              unloadMuxOut[17] = fifoOut[38][16][w-1];
              unloadMuxOut[18] = fifoOut[39][16][w-1];
              unloadMuxOut[19] = fifoOut[40][16][w-1];
              unloadMuxOut[20] = fifoOut[41][16][w-1];
              unloadMuxOut[21] = fifoOut[42][16][w-1];
              unloadMuxOut[22] = fifoOut[43][16][w-1];
              unloadMuxOut[23] = fifoOut[44][16][w-1];
              unloadMuxOut[24] = fifoOut[45][16][w-1];
              unloadMuxOut[25] = fifoOut[46][16][w-1];
              unloadMuxOut[26] = fifoOut[47][16][w-1];
              unloadMuxOut[27] = fifoOut[48][16][w-1];
              unloadMuxOut[28] = fifoOut[49][16][w-1];
              unloadMuxOut[29] = fifoOut[50][16][w-1];
              unloadMuxOut[30] = fifoOut[51][16][w-1];
              unloadMuxOut[31] = fifoOut[26][15][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[27][16][w-1];
              unloadMuxOut[1] = fifoOut[28][16][w-1];
              unloadMuxOut[2] = fifoOut[29][16][w-1];
              unloadMuxOut[3] = fifoOut[30][16][w-1];
              unloadMuxOut[4] = fifoOut[31][16][w-1];
              unloadMuxOut[5] = fifoOut[32][16][w-1];
              unloadMuxOut[6] = fifoOut[33][16][w-1];
              unloadMuxOut[7] = fifoOut[34][16][w-1];
              unloadMuxOut[8] = fifoOut[35][16][w-1];
              unloadMuxOut[9] = fifoOut[36][16][w-1];
              unloadMuxOut[10] = fifoOut[37][16][w-1];
              unloadMuxOut[11] = fifoOut[38][16][w-1];
              unloadMuxOut[12] = fifoOut[39][16][w-1];
              unloadMuxOut[13] = fifoOut[40][16][w-1];
              unloadMuxOut[14] = fifoOut[41][16][w-1];
              unloadMuxOut[15] = fifoOut[42][16][w-1];
              unloadMuxOut[16] = fifoOut[43][16][w-1];
              unloadMuxOut[17] = fifoOut[44][16][w-1];
              unloadMuxOut[18] = fifoOut[45][16][w-1];
              unloadMuxOut[19] = fifoOut[46][16][w-1];
              unloadMuxOut[20] = fifoOut[47][16][w-1];
              unloadMuxOut[21] = fifoOut[48][16][w-1];
              unloadMuxOut[22] = fifoOut[49][16][w-1];
              unloadMuxOut[23] = fifoOut[50][16][w-1];
              unloadMuxOut[24] = fifoOut[51][16][w-1];
              unloadMuxOut[25] = fifoOut[26][15][w-1];
              unloadMuxOut[26] = fifoOut[27][15][w-1];
              unloadMuxOut[27] = fifoOut[28][15][w-1];
              unloadMuxOut[28] = fifoOut[29][15][w-1];
              unloadMuxOut[29] = fifoOut[30][15][w-1];
              unloadMuxOut[30] = fifoOut[31][15][w-1];
              unloadMuxOut[31] = fifoOut[32][15][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[33][16][w-1];
              unloadMuxOut[1] = fifoOut[34][16][w-1];
              unloadMuxOut[2] = fifoOut[35][16][w-1];
              unloadMuxOut[3] = fifoOut[36][16][w-1];
              unloadMuxOut[4] = fifoOut[37][16][w-1];
              unloadMuxOut[5] = fifoOut[38][16][w-1];
              unloadMuxOut[6] = fifoOut[39][16][w-1];
              unloadMuxOut[7] = fifoOut[40][16][w-1];
              unloadMuxOut[8] = fifoOut[41][16][w-1];
              unloadMuxOut[9] = fifoOut[42][16][w-1];
              unloadMuxOut[10] = fifoOut[43][16][w-1];
              unloadMuxOut[11] = fifoOut[44][16][w-1];
              unloadMuxOut[12] = fifoOut[45][16][w-1];
              unloadMuxOut[13] = fifoOut[46][16][w-1];
              unloadMuxOut[14] = fifoOut[47][16][w-1];
              unloadMuxOut[15] = fifoOut[48][16][w-1];
              unloadMuxOut[16] = fifoOut[49][16][w-1];
              unloadMuxOut[17] = fifoOut[50][16][w-1];
              unloadMuxOut[18] = fifoOut[51][16][w-1];
              unloadMuxOut[19] = fifoOut[26][15][w-1];
              unloadMuxOut[20] = fifoOut[27][15][w-1];
              unloadMuxOut[21] = fifoOut[28][15][w-1];
              unloadMuxOut[22] = fifoOut[29][15][w-1];
              unloadMuxOut[23] = fifoOut[30][15][w-1];
              unloadMuxOut[24] = fifoOut[31][15][w-1];
              unloadMuxOut[25] = fifoOut[32][15][w-1];
              unloadMuxOut[26] = fifoOut[33][15][w-1];
              unloadMuxOut[27] = fifoOut[34][15][w-1];
              unloadMuxOut[28] = fifoOut[35][15][w-1];
              unloadMuxOut[29] = fifoOut[36][15][w-1];
              unloadMuxOut[30] = fifoOut[37][15][w-1];
              unloadMuxOut[31] = fifoOut[38][15][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[39][16][w-1];
              unloadMuxOut[1] = fifoOut[40][16][w-1];
              unloadMuxOut[2] = fifoOut[41][16][w-1];
              unloadMuxOut[3] = fifoOut[42][16][w-1];
              unloadMuxOut[4] = fifoOut[43][16][w-1];
              unloadMuxOut[5] = fifoOut[44][16][w-1];
              unloadMuxOut[6] = fifoOut[45][16][w-1];
              unloadMuxOut[7] = fifoOut[46][16][w-1];
              unloadMuxOut[8] = fifoOut[47][16][w-1];
              unloadMuxOut[9] = fifoOut[48][16][w-1];
              unloadMuxOut[10] = fifoOut[49][16][w-1];
              unloadMuxOut[11] = fifoOut[50][16][w-1];
              unloadMuxOut[12] = fifoOut[51][16][w-1];
              unloadMuxOut[13] = fifoOut[26][15][w-1];
              unloadMuxOut[14] = fifoOut[27][15][w-1];
              unloadMuxOut[15] = fifoOut[28][15][w-1];
              unloadMuxOut[16] = fifoOut[29][15][w-1];
              unloadMuxOut[17] = fifoOut[30][15][w-1];
              unloadMuxOut[18] = fifoOut[31][15][w-1];
              unloadMuxOut[19] = fifoOut[32][15][w-1];
              unloadMuxOut[20] = fifoOut[33][15][w-1];
              unloadMuxOut[21] = fifoOut[34][15][w-1];
              unloadMuxOut[22] = fifoOut[35][15][w-1];
              unloadMuxOut[23] = fifoOut[36][15][w-1];
              unloadMuxOut[24] = fifoOut[37][15][w-1];
              unloadMuxOut[25] = fifoOut[38][15][w-1];
              unloadMuxOut[26] = fifoOut[39][15][w-1];
              unloadMuxOut[27] = fifoOut[40][15][w-1];
              unloadMuxOut[28] = fifoOut[41][15][w-1];
              unloadMuxOut[29] = fifoOut[42][15][w-1];
              unloadMuxOut[30] = fifoOut[43][15][w-1];
              unloadMuxOut[31] = fifoOut[44][15][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[45][16][w-1];
              unloadMuxOut[1] = fifoOut[46][16][w-1];
              unloadMuxOut[2] = fifoOut[47][16][w-1];
              unloadMuxOut[3] = fifoOut[48][16][w-1];
              unloadMuxOut[4] = fifoOut[49][16][w-1];
              unloadMuxOut[5] = fifoOut[50][16][w-1];
              unloadMuxOut[6] = fifoOut[51][16][w-1];
              unloadMuxOut[7] = fifoOut[26][15][w-1];
              unloadMuxOut[8] = fifoOut[27][15][w-1];
              unloadMuxOut[9] = fifoOut[28][15][w-1];
              unloadMuxOut[10] = fifoOut[29][15][w-1];
              unloadMuxOut[11] = fifoOut[30][15][w-1];
              unloadMuxOut[12] = fifoOut[31][15][w-1];
              unloadMuxOut[13] = fifoOut[32][15][w-1];
              unloadMuxOut[14] = fifoOut[33][15][w-1];
              unloadMuxOut[15] = fifoOut[34][15][w-1];
              unloadMuxOut[16] = fifoOut[35][15][w-1];
              unloadMuxOut[17] = fifoOut[36][15][w-1];
              unloadMuxOut[18] = fifoOut[37][15][w-1];
              unloadMuxOut[19] = fifoOut[38][15][w-1];
              unloadMuxOut[20] = fifoOut[39][15][w-1];
              unloadMuxOut[21] = fifoOut[40][15][w-1];
              unloadMuxOut[22] = fifoOut[41][15][w-1];
              unloadMuxOut[23] = fifoOut[42][15][w-1];
              unloadMuxOut[24] = fifoOut[43][15][w-1];
              unloadMuxOut[25] = fifoOut[44][15][w-1];
              unloadMuxOut[26] = fifoOut[45][15][w-1];
              unloadMuxOut[27] = fifoOut[46][15][w-1];
              unloadMuxOut[28] = fifoOut[47][15][w-1];
              unloadMuxOut[29] = fifoOut[48][15][w-1];
              unloadMuxOut[30] = fifoOut[49][15][w-1];
              unloadMuxOut[31] = fifoOut[50][15][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[51][16][w-1];
              unloadMuxOut[1] = fifoOut[26][15][w-1];
              unloadMuxOut[2] = fifoOut[27][15][w-1];
              unloadMuxOut[3] = fifoOut[28][15][w-1];
              unloadMuxOut[4] = fifoOut[29][15][w-1];
              unloadMuxOut[5] = fifoOut[30][15][w-1];
              unloadMuxOut[6] = fifoOut[31][15][w-1];
              unloadMuxOut[7] = fifoOut[32][15][w-1];
              unloadMuxOut[8] = fifoOut[33][15][w-1];
              unloadMuxOut[9] = fifoOut[34][15][w-1];
              unloadMuxOut[10] = fifoOut[35][15][w-1];
              unloadMuxOut[11] = fifoOut[36][15][w-1];
              unloadMuxOut[12] = fifoOut[37][15][w-1];
              unloadMuxOut[13] = fifoOut[38][15][w-1];
              unloadMuxOut[14] = fifoOut[39][15][w-1];
              unloadMuxOut[15] = fifoOut[40][15][w-1];
              unloadMuxOut[16] = fifoOut[41][15][w-1];
              unloadMuxOut[17] = fifoOut[42][15][w-1];
              unloadMuxOut[18] = fifoOut[43][15][w-1];
              unloadMuxOut[19] = fifoOut[44][15][w-1];
              unloadMuxOut[20] = fifoOut[45][15][w-1];
              unloadMuxOut[21] = fifoOut[46][15][w-1];
              unloadMuxOut[22] = fifoOut[47][15][w-1];
              unloadMuxOut[23] = fifoOut[48][15][w-1];
              unloadMuxOut[24] = fifoOut[49][15][w-1];
              unloadMuxOut[25] = fifoOut[50][15][w-1];
              unloadMuxOut[26] = fifoOut[51][15][w-1];
              unloadMuxOut[27] = fifoOut[26][14][w-1];
              unloadMuxOut[28] = fifoOut[27][14][w-1];
              unloadMuxOut[29] = fifoOut[28][14][w-1];
              unloadMuxOut[30] = fifoOut[29][14][w-1];
              unloadMuxOut[31] = fifoOut[30][14][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[31][15][w-1];
              unloadMuxOut[1] = fifoOut[32][15][w-1];
              unloadMuxOut[2] = fifoOut[33][15][w-1];
              unloadMuxOut[3] = fifoOut[34][15][w-1];
              unloadMuxOut[4] = fifoOut[35][15][w-1];
              unloadMuxOut[5] = fifoOut[36][15][w-1];
              unloadMuxOut[6] = fifoOut[37][15][w-1];
              unloadMuxOut[7] = fifoOut[38][15][w-1];
              unloadMuxOut[8] = fifoOut[39][15][w-1];
              unloadMuxOut[9] = fifoOut[40][15][w-1];
              unloadMuxOut[10] = fifoOut[41][15][w-1];
              unloadMuxOut[11] = fifoOut[42][15][w-1];
              unloadMuxOut[12] = fifoOut[43][15][w-1];
              unloadMuxOut[13] = fifoOut[44][15][w-1];
              unloadMuxOut[14] = fifoOut[45][15][w-1];
              unloadMuxOut[15] = fifoOut[46][15][w-1];
              unloadMuxOut[16] = fifoOut[47][15][w-1];
              unloadMuxOut[17] = fifoOut[48][15][w-1];
              unloadMuxOut[18] = fifoOut[49][15][w-1];
              unloadMuxOut[19] = fifoOut[50][15][w-1];
              unloadMuxOut[20] = fifoOut[51][15][w-1];
              unloadMuxOut[21] = fifoOut[26][14][w-1];
              unloadMuxOut[22] = fifoOut[27][14][w-1];
              unloadMuxOut[23] = fifoOut[28][14][w-1];
              unloadMuxOut[24] = fifoOut[29][14][w-1];
              unloadMuxOut[25] = fifoOut[30][14][w-1];
              unloadMuxOut[26] = fifoOut[31][14][w-1];
              unloadMuxOut[27] = fifoOut[32][14][w-1];
              unloadMuxOut[28] = fifoOut[33][14][w-1];
              unloadMuxOut[29] = fifoOut[34][14][w-1];
              unloadMuxOut[30] = fifoOut[35][14][w-1];
              unloadMuxOut[31] = fifoOut[36][14][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[37][15][w-1];
              unloadMuxOut[1] = fifoOut[38][15][w-1];
              unloadMuxOut[2] = fifoOut[39][15][w-1];
              unloadMuxOut[3] = fifoOut[40][15][w-1];
              unloadMuxOut[4] = fifoOut[41][15][w-1];
              unloadMuxOut[5] = fifoOut[42][15][w-1];
              unloadMuxOut[6] = fifoOut[43][15][w-1];
              unloadMuxOut[7] = fifoOut[44][15][w-1];
              unloadMuxOut[8] = fifoOut[45][15][w-1];
              unloadMuxOut[9] = fifoOut[46][15][w-1];
              unloadMuxOut[10] = fifoOut[47][15][w-1];
              unloadMuxOut[11] = fifoOut[48][15][w-1];
              unloadMuxOut[12] = fifoOut[49][15][w-1];
              unloadMuxOut[13] = fifoOut[50][15][w-1];
              unloadMuxOut[14] = fifoOut[51][15][w-1];
              unloadMuxOut[15] = fifoOut[26][14][w-1];
              unloadMuxOut[16] = fifoOut[27][14][w-1];
              unloadMuxOut[17] = fifoOut[28][14][w-1];
              unloadMuxOut[18] = fifoOut[29][14][w-1];
              unloadMuxOut[19] = fifoOut[30][14][w-1];
              unloadMuxOut[20] = fifoOut[31][14][w-1];
              unloadMuxOut[21] = fifoOut[32][14][w-1];
              unloadMuxOut[22] = fifoOut[33][14][w-1];
              unloadMuxOut[23] = fifoOut[34][14][w-1];
              unloadMuxOut[24] = fifoOut[35][14][w-1];
              unloadMuxOut[25] = fifoOut[36][14][w-1];
              unloadMuxOut[26] = fifoOut[37][14][w-1];
              unloadMuxOut[27] = fifoOut[38][14][w-1];
              unloadMuxOut[28] = fifoOut[39][14][w-1];
              unloadMuxOut[29] = fifoOut[40][14][w-1];
              unloadMuxOut[30] = fifoOut[41][14][w-1];
              unloadMuxOut[31] = fifoOut[42][14][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[43][15][w-1];
              unloadMuxOut[1] = fifoOut[44][15][w-1];
              unloadMuxOut[2] = fifoOut[45][15][w-1];
              unloadMuxOut[3] = fifoOut[46][15][w-1];
              unloadMuxOut[4] = fifoOut[47][15][w-1];
              unloadMuxOut[5] = fifoOut[48][15][w-1];
              unloadMuxOut[6] = fifoOut[49][15][w-1];
              unloadMuxOut[7] = fifoOut[50][15][w-1];
              unloadMuxOut[8] = fifoOut[51][15][w-1];
              unloadMuxOut[9] = fifoOut[26][14][w-1];
              unloadMuxOut[10] = fifoOut[27][14][w-1];
              unloadMuxOut[11] = fifoOut[28][14][w-1];
              unloadMuxOut[12] = fifoOut[29][14][w-1];
              unloadMuxOut[13] = fifoOut[30][14][w-1];
              unloadMuxOut[14] = fifoOut[31][14][w-1];
              unloadMuxOut[15] = fifoOut[32][14][w-1];
              unloadMuxOut[16] = fifoOut[33][14][w-1];
              unloadMuxOut[17] = fifoOut[34][14][w-1];
              unloadMuxOut[18] = fifoOut[35][14][w-1];
              unloadMuxOut[19] = fifoOut[36][14][w-1];
              unloadMuxOut[20] = fifoOut[37][14][w-1];
              unloadMuxOut[21] = fifoOut[38][14][w-1];
              unloadMuxOut[22] = fifoOut[39][14][w-1];
              unloadMuxOut[23] = fifoOut[40][14][w-1];
              unloadMuxOut[24] = fifoOut[41][14][w-1];
              unloadMuxOut[25] = fifoOut[42][14][w-1];
              unloadMuxOut[26] = fifoOut[19][11][w-1];
              unloadMuxOut[27] = fifoOut[20][11][w-1];
              unloadMuxOut[28] = fifoOut[21][11][w-1];
              unloadMuxOut[29] = fifoOut[22][11][w-1];
              unloadMuxOut[30] = fifoOut[23][11][w-1];
              unloadMuxOut[31] = fifoOut[24][11][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[25][12][w-1];
              unloadMuxOut[1] = fifoOut[0][11][w-1];
              unloadMuxOut[2] = fifoOut[1][11][w-1];
              unloadMuxOut[3] = fifoOut[2][11][w-1];
              unloadMuxOut[4] = fifoOut[3][11][w-1];
              unloadMuxOut[5] = fifoOut[4][11][w-1];
              unloadMuxOut[6] = fifoOut[5][11][w-1];
              unloadMuxOut[7] = fifoOut[6][11][w-1];
              unloadMuxOut[8] = fifoOut[7][11][w-1];
              unloadMuxOut[9] = fifoOut[8][11][w-1];
              unloadMuxOut[10] = fifoOut[9][11][w-1];
              unloadMuxOut[11] = fifoOut[10][11][w-1];
              unloadMuxOut[12] = fifoOut[11][11][w-1];
              unloadMuxOut[13] = fifoOut[12][11][w-1];
              unloadMuxOut[14] = fifoOut[13][11][w-1];
              unloadMuxOut[15] = fifoOut[14][11][w-1];
              unloadMuxOut[16] = fifoOut[15][11][w-1];
              unloadMuxOut[17] = fifoOut[16][11][w-1];
              unloadMuxOut[18] = fifoOut[17][11][w-1];
              unloadMuxOut[19] = fifoOut[18][11][w-1];
              unloadMuxOut[20] = fifoOut[19][11][w-1];
              unloadMuxOut[21] = fifoOut[20][11][w-1];
              unloadMuxOut[22] = fifoOut[21][11][w-1];
              unloadMuxOut[23] = fifoOut[22][11][w-1];
              unloadMuxOut[24] = fifoOut[23][11][w-1];
              unloadMuxOut[25] = fifoOut[24][11][w-1];
              unloadMuxOut[26] = fifoOut[25][11][w-1];
              unloadMuxOut[27] = fifoOut[0][10][w-1];
              unloadMuxOut[28] = fifoOut[1][10][w-1];
              unloadMuxOut[29] = fifoOut[2][10][w-1];
              unloadMuxOut[30] = fifoOut[3][10][w-1];
              unloadMuxOut[31] = fifoOut[4][10][w-1];
       end
       16: begin
              unloadMuxOut[0] = fifoOut[5][11][w-1];
              unloadMuxOut[1] = fifoOut[6][11][w-1];
              unloadMuxOut[2] = fifoOut[7][11][w-1];
              unloadMuxOut[3] = fifoOut[8][11][w-1];
              unloadMuxOut[4] = fifoOut[9][11][w-1];
              unloadMuxOut[5] = fifoOut[10][11][w-1];
              unloadMuxOut[6] = fifoOut[11][11][w-1];
              unloadMuxOut[7] = fifoOut[12][11][w-1];
              unloadMuxOut[8] = fifoOut[13][11][w-1];
              unloadMuxOut[9] = fifoOut[14][11][w-1];
              unloadMuxOut[10] = fifoOut[15][11][w-1];
              unloadMuxOut[11] = fifoOut[16][11][w-1];
              unloadMuxOut[12] = fifoOut[17][11][w-1];
              unloadMuxOut[13] = fifoOut[18][11][w-1];
              unloadMuxOut[14] = fifoOut[19][11][w-1];
              unloadMuxOut[15] = fifoOut[20][11][w-1];
              unloadMuxOut[16] = fifoOut[21][11][w-1];
              unloadMuxOut[17] = fifoOut[22][11][w-1];
              unloadMuxOut[18] = fifoOut[23][11][w-1];
              unloadMuxOut[19] = fifoOut[24][11][w-1];
              unloadMuxOut[20] = fifoOut[25][11][w-1];
              unloadMuxOut[21] = fifoOut[0][10][w-1];
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0; 
             end
       end
    endcase //unload case end
    case(iteration_0_indicator)
       0: begin
         case(rd_address_case)
         0: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[43][4];
              muxOutConnector[45] = fifoOut[44][4];
              muxOutConnector[46] = fifoOut[45][4];
              muxOutConnector[47] = fifoOut[46][4];
              muxOutConnector[48] = fifoOut[47][4];
              muxOutConnector[49] = fifoOut[48][4];
              muxOutConnector[50] = fifoOut[49][4];
              muxOutConnector[51] = fifoOut[50][4];
         end
         1: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[43][15];
              muxOutConnector[9] = fifoOut[44][15];
              muxOutConnector[10] = fifoOut[45][15];
              muxOutConnector[11] = fifoOut[46][15];
              muxOutConnector[12] = fifoOut[47][15];
              muxOutConnector[13] = fifoOut[48][15];
              muxOutConnector[14] = fifoOut[49][15];
              muxOutConnector[15] = fifoOut[50][15];
              muxOutConnector[16] = fifoOut[51][15];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[43][4];
              muxOutConnector[45] = fifoOut[44][4];
              muxOutConnector[46] = fifoOut[45][4];
              muxOutConnector[47] = fifoOut[46][4];
              muxOutConnector[48] = fifoOut[47][4];
              muxOutConnector[49] = fifoOut[48][4];
              muxOutConnector[50] = fifoOut[49][4];
              muxOutConnector[51] = fifoOut[50][4];
         end
         2: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[43][15];
              muxOutConnector[9] = fifoOut[44][15];
              muxOutConnector[10] = fifoOut[45][15];
              muxOutConnector[11] = fifoOut[46][15];
              muxOutConnector[12] = fifoOut[47][15];
              muxOutConnector[13] = fifoOut[48][15];
              muxOutConnector[14] = fifoOut[49][15];
              muxOutConnector[15] = fifoOut[50][15];
              muxOutConnector[16] = fifoOut[51][15];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[43][4];
              muxOutConnector[45] = fifoOut[44][4];
              muxOutConnector[46] = fifoOut[45][4];
              muxOutConnector[47] = fifoOut[46][4];
              muxOutConnector[48] = fifoOut[47][4];
              muxOutConnector[49] = fifoOut[48][4];
              muxOutConnector[50] = fifoOut[49][4];
              muxOutConnector[51] = fifoOut[50][4];
         end
         3: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[43][15];
              muxOutConnector[9] = fifoOut[44][15];
              muxOutConnector[10] = fifoOut[45][15];
              muxOutConnector[11] = fifoOut[46][15];
              muxOutConnector[12] = fifoOut[47][15];
              muxOutConnector[13] = fifoOut[48][15];
              muxOutConnector[14] = fifoOut[49][15];
              muxOutConnector[15] = fifoOut[50][15];
              muxOutConnector[16] = fifoOut[51][15];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[43][4];
              muxOutConnector[45] = fifoOut[44][4];
              muxOutConnector[46] = fifoOut[45][4];
              muxOutConnector[47] = fifoOut[46][4];
              muxOutConnector[48] = fifoOut[47][4];
              muxOutConnector[49] = fifoOut[48][4];
              muxOutConnector[50] = fifoOut[49][4];
              muxOutConnector[51] = fifoOut[50][4];
         end
         4: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[43][15];
              muxOutConnector[9] = fifoOut[44][15];
              muxOutConnector[10] = fifoOut[45][15];
              muxOutConnector[11] = fifoOut[46][15];
              muxOutConnector[12] = fifoOut[47][15];
              muxOutConnector[13] = fifoOut[48][15];
              muxOutConnector[14] = fifoOut[49][15];
              muxOutConnector[15] = fifoOut[50][15];
              muxOutConnector[16] = fifoOut[51][15];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[19][1];
              muxOutConnector[45] = fifoOut[20][1];
              muxOutConnector[46] = fifoOut[21][1];
              muxOutConnector[47] = fifoOut[22][1];
              muxOutConnector[48] = fifoOut[23][1];
              muxOutConnector[49] = fifoOut[24][1];
              muxOutConnector[50] = fifoOut[25][1];
              muxOutConnector[51] = fifoOut[0][0];
         end
         5: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[43][15];
              muxOutConnector[9] = fifoOut[44][15];
              muxOutConnector[10] = fifoOut[45][15];
              muxOutConnector[11] = fifoOut[46][15];
              muxOutConnector[12] = fifoOut[47][15];
              muxOutConnector[13] = fifoOut[48][15];
              muxOutConnector[14] = fifoOut[49][15];
              muxOutConnector[15] = fifoOut[50][15];
              muxOutConnector[16] = fifoOut[51][15];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][1];
              muxOutConnector[27] = fifoOut[2][1];
              muxOutConnector[28] = fifoOut[3][1];
              muxOutConnector[29] = fifoOut[4][1];
              muxOutConnector[30] = fifoOut[5][1];
              muxOutConnector[31] = fifoOut[6][1];
              muxOutConnector[32] = fifoOut[7][1];
              muxOutConnector[33] = fifoOut[8][1];
              muxOutConnector[34] = fifoOut[9][1];
              muxOutConnector[35] = fifoOut[10][1];
              muxOutConnector[36] = fifoOut[11][1];
              muxOutConnector[37] = fifoOut[12][1];
              muxOutConnector[38] = fifoOut[13][1];
              muxOutConnector[39] = fifoOut[14][1];
              muxOutConnector[40] = fifoOut[15][1];
              muxOutConnector[41] = fifoOut[16][1];
              muxOutConnector[42] = fifoOut[17][1];
              muxOutConnector[43] = fifoOut[18][1];
              muxOutConnector[44] = fifoOut[19][1];
              muxOutConnector[45] = fifoOut[20][1];
              muxOutConnector[46] = fifoOut[21][1];
              muxOutConnector[47] = fifoOut[22][1];
              muxOutConnector[48] = fifoOut[23][1];
              muxOutConnector[49] = fifoOut[24][1];
              muxOutConnector[50] = fifoOut[25][1];
              muxOutConnector[51] = fifoOut[0][0];
         end
         6: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[43][15];
              muxOutConnector[9] = fifoOut[44][15];
              muxOutConnector[10] = fifoOut[45][15];
              muxOutConnector[11] = fifoOut[46][15];
              muxOutConnector[12] = fifoOut[47][15];
              muxOutConnector[13] = fifoOut[48][15];
              muxOutConnector[14] = fifoOut[49][15];
              muxOutConnector[15] = fifoOut[50][15];
              muxOutConnector[16] = fifoOut[51][15];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][1];
              muxOutConnector[27] = fifoOut[2][1];
              muxOutConnector[28] = fifoOut[3][1];
              muxOutConnector[29] = fifoOut[4][1];
              muxOutConnector[30] = fifoOut[5][1];
              muxOutConnector[31] = fifoOut[6][1];
              muxOutConnector[32] = fifoOut[7][1];
              muxOutConnector[33] = fifoOut[8][1];
              muxOutConnector[34] = fifoOut[9][1];
              muxOutConnector[35] = fifoOut[10][1];
              muxOutConnector[36] = fifoOut[11][1];
              muxOutConnector[37] = fifoOut[12][1];
              muxOutConnector[38] = fifoOut[13][1];
              muxOutConnector[39] = fifoOut[14][1];
              muxOutConnector[40] = fifoOut[15][1];
              muxOutConnector[41] = fifoOut[16][1];
              muxOutConnector[42] = fifoOut[17][1];
              muxOutConnector[43] = fifoOut[18][1];
              muxOutConnector[44] = fifoOut[19][1];
              muxOutConnector[45] = fifoOut[20][1];
              muxOutConnector[46] = fifoOut[21][1];
              muxOutConnector[47] = fifoOut[22][1];
              muxOutConnector[48] = fifoOut[23][1];
              muxOutConnector[49] = fifoOut[24][1];
              muxOutConnector[50] = fifoOut[25][1];
              muxOutConnector[51] = fifoOut[0][0];
         end
         7: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[43][15];
              muxOutConnector[9] = fifoOut[44][15];
              muxOutConnector[10] = fifoOut[45][15];
              muxOutConnector[11] = fifoOut[46][15];
              muxOutConnector[12] = fifoOut[47][15];
              muxOutConnector[13] = fifoOut[48][15];
              muxOutConnector[14] = fifoOut[49][15];
              muxOutConnector[15] = fifoOut[50][15];
              muxOutConnector[16] = fifoOut[51][15];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][1];
              muxOutConnector[27] = fifoOut[2][1];
              muxOutConnector[28] = fifoOut[3][1];
              muxOutConnector[29] = fifoOut[4][1];
              muxOutConnector[30] = fifoOut[5][1];
              muxOutConnector[31] = fifoOut[6][1];
              muxOutConnector[32] = fifoOut[7][1];
              muxOutConnector[33] = fifoOut[8][1];
              muxOutConnector[34] = fifoOut[9][1];
              muxOutConnector[35] = fifoOut[10][1];
              muxOutConnector[36] = fifoOut[11][1];
              muxOutConnector[37] = fifoOut[12][1];
              muxOutConnector[38] = fifoOut[13][1];
              muxOutConnector[39] = fifoOut[14][1];
              muxOutConnector[40] = fifoOut[15][1];
              muxOutConnector[41] = fifoOut[16][1];
              muxOutConnector[42] = fifoOut[17][1];
              muxOutConnector[43] = fifoOut[18][1];
              muxOutConnector[44] = fifoOut[19][1];
              muxOutConnector[45] = fifoOut[20][1];
              muxOutConnector[46] = fifoOut[21][1];
              muxOutConnector[47] = fifoOut[22][1];
              muxOutConnector[48] = fifoOut[23][1];
              muxOutConnector[49] = fifoOut[24][1];
              muxOutConnector[50] = fifoOut[25][1];
              muxOutConnector[51] = fifoOut[0][0];
         end
         8: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[43][15];
              muxOutConnector[9] = fifoOut[44][15];
              muxOutConnector[10] = fifoOut[45][15];
              muxOutConnector[11] = fifoOut[46][15];
              muxOutConnector[12] = fifoOut[47][15];
              muxOutConnector[13] = fifoOut[48][15];
              muxOutConnector[14] = fifoOut[49][15];
              muxOutConnector[15] = fifoOut[50][15];
              muxOutConnector[16] = fifoOut[51][15];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][1];
              muxOutConnector[27] = fifoOut[2][1];
              muxOutConnector[28] = fifoOut[3][1];
              muxOutConnector[29] = fifoOut[4][1];
              muxOutConnector[30] = fifoOut[5][1];
              muxOutConnector[31] = fifoOut[6][1];
              muxOutConnector[32] = fifoOut[7][1];
              muxOutConnector[33] = fifoOut[8][1];
              muxOutConnector[34] = fifoOut[9][1];
              muxOutConnector[35] = fifoOut[10][1];
              muxOutConnector[36] = fifoOut[11][1];
              muxOutConnector[37] = fifoOut[12][1];
              muxOutConnector[38] = fifoOut[13][1];
              muxOutConnector[39] = fifoOut[14][1];
              muxOutConnector[40] = fifoOut[15][1];
              muxOutConnector[41] = fifoOut[16][1];
              muxOutConnector[42] = fifoOut[17][1];
              muxOutConnector[43] = fifoOut[18][1];
              muxOutConnector[44] = fifoOut[19][1];
              muxOutConnector[45] = fifoOut[20][1];
              muxOutConnector[46] = fifoOut[21][1];
              muxOutConnector[47] = fifoOut[22][1];
              muxOutConnector[48] = fifoOut[23][1];
              muxOutConnector[49] = fifoOut[24][1];
              muxOutConnector[50] = fifoOut[25][1];
              muxOutConnector[51] = fifoOut[0][0];
         end
         9: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[43][15];
              muxOutConnector[9] = fifoOut[44][15];
              muxOutConnector[10] = fifoOut[45][15];
              muxOutConnector[11] = fifoOut[46][15];
              muxOutConnector[12] = fifoOut[47][15];
              muxOutConnector[13] = fifoOut[48][15];
              muxOutConnector[14] = fifoOut[49][15];
              muxOutConnector[15] = fifoOut[50][15];
              muxOutConnector[16] = fifoOut[51][15];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][1];
              muxOutConnector[27] = fifoOut[2][1];
              muxOutConnector[28] = fifoOut[3][1];
              muxOutConnector[29] = fifoOut[4][1];
              muxOutConnector[30] = fifoOut[5][1];
              muxOutConnector[31] = fifoOut[6][1];
              muxOutConnector[32] = fifoOut[7][1];
              muxOutConnector[33] = fifoOut[8][1];
              muxOutConnector[34] = fifoOut[9][1];
              muxOutConnector[35] = fifoOut[10][1];
              muxOutConnector[36] = fifoOut[11][1];
              muxOutConnector[37] = fifoOut[12][1];
              muxOutConnector[38] = fifoOut[13][1];
              muxOutConnector[39] = fifoOut[14][1];
              muxOutConnector[40] = fifoOut[15][1];
              muxOutConnector[41] = fifoOut[16][1];
              muxOutConnector[42] = fifoOut[17][1];
              muxOutConnector[43] = fifoOut[18][1];
              muxOutConnector[44] = fifoOut[26][6];
              muxOutConnector[45] = fifoOut[27][6];
              muxOutConnector[46] = fifoOut[28][6];
              muxOutConnector[47] = fifoOut[29][6];
              muxOutConnector[48] = fifoOut[30][6];
              muxOutConnector[49] = fifoOut[31][6];
              muxOutConnector[50] = fifoOut[32][6];
              muxOutConnector[51] = fifoOut[33][6];
         end
         10: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[43][15];
              muxOutConnector[9] = fifoOut[44][15];
              muxOutConnector[10] = fifoOut[45][15];
              muxOutConnector[11] = fifoOut[46][15];
              muxOutConnector[12] = fifoOut[47][15];
              muxOutConnector[13] = fifoOut[48][15];
              muxOutConnector[14] = fifoOut[49][15];
              muxOutConnector[15] = fifoOut[50][15];
              muxOutConnector[16] = fifoOut[51][15];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][7];
              muxOutConnector[27] = fifoOut[35][7];
              muxOutConnector[28] = fifoOut[36][7];
              muxOutConnector[29] = fifoOut[37][7];
              muxOutConnector[30] = fifoOut[38][7];
              muxOutConnector[31] = fifoOut[39][7];
              muxOutConnector[32] = fifoOut[40][7];
              muxOutConnector[33] = fifoOut[41][7];
              muxOutConnector[34] = fifoOut[42][7];
              muxOutConnector[35] = fifoOut[43][7];
              muxOutConnector[36] = fifoOut[44][7];
              muxOutConnector[37] = fifoOut[45][7];
              muxOutConnector[38] = fifoOut[46][7];
              muxOutConnector[39] = fifoOut[47][7];
              muxOutConnector[40] = fifoOut[48][7];
              muxOutConnector[41] = fifoOut[49][7];
              muxOutConnector[42] = fifoOut[50][7];
              muxOutConnector[43] = fifoOut[51][7];
              muxOutConnector[44] = fifoOut[26][6];
              muxOutConnector[45] = fifoOut[27][6];
              muxOutConnector[46] = fifoOut[28][6];
              muxOutConnector[47] = fifoOut[29][6];
              muxOutConnector[48] = fifoOut[30][6];
              muxOutConnector[49] = fifoOut[31][6];
              muxOutConnector[50] = fifoOut[32][6];
              muxOutConnector[51] = fifoOut[33][6];
         end
         11: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[43][15];
              muxOutConnector[9] = fifoOut[44][15];
              muxOutConnector[10] = fifoOut[45][15];
              muxOutConnector[11] = fifoOut[46][15];
              muxOutConnector[12] = fifoOut[47][15];
              muxOutConnector[13] = fifoOut[48][15];
              muxOutConnector[14] = fifoOut[49][15];
              muxOutConnector[15] = fifoOut[50][15];
              muxOutConnector[16] = fifoOut[51][15];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][7];
              muxOutConnector[27] = fifoOut[35][7];
              muxOutConnector[28] = fifoOut[36][7];
              muxOutConnector[29] = fifoOut[37][7];
              muxOutConnector[30] = fifoOut[38][7];
              muxOutConnector[31] = fifoOut[39][7];
              muxOutConnector[32] = fifoOut[40][7];
              muxOutConnector[33] = fifoOut[41][7];
              muxOutConnector[34] = fifoOut[42][7];
              muxOutConnector[35] = fifoOut[43][7];
              muxOutConnector[36] = fifoOut[44][7];
              muxOutConnector[37] = fifoOut[45][7];
              muxOutConnector[38] = fifoOut[46][7];
              muxOutConnector[39] = fifoOut[47][7];
              muxOutConnector[40] = fifoOut[48][7];
              muxOutConnector[41] = fifoOut[49][7];
              muxOutConnector[42] = fifoOut[50][7];
              muxOutConnector[43] = fifoOut[51][7];
              muxOutConnector[44] = fifoOut[26][6];
              muxOutConnector[45] = fifoOut[27][6];
              muxOutConnector[46] = fifoOut[28][6];
              muxOutConnector[47] = fifoOut[29][6];
              muxOutConnector[48] = fifoOut[30][6];
              muxOutConnector[49] = fifoOut[31][6];
              muxOutConnector[50] = fifoOut[32][6];
              muxOutConnector[51] = fifoOut[33][6];
         end
         12: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[43][15];
              muxOutConnector[9] = fifoOut[44][15];
              muxOutConnector[10] = fifoOut[45][15];
              muxOutConnector[11] = fifoOut[46][15];
              muxOutConnector[12] = fifoOut[47][15];
              muxOutConnector[13] = fifoOut[48][15];
              muxOutConnector[14] = fifoOut[49][15];
              muxOutConnector[15] = fifoOut[50][15];
              muxOutConnector[16] = fifoOut[51][15];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][7];
              muxOutConnector[27] = fifoOut[35][7];
              muxOutConnector[28] = fifoOut[36][7];
              muxOutConnector[29] = fifoOut[37][7];
              muxOutConnector[30] = fifoOut[38][7];
              muxOutConnector[31] = fifoOut[39][7];
              muxOutConnector[32] = fifoOut[40][7];
              muxOutConnector[33] = fifoOut[41][7];
              muxOutConnector[34] = fifoOut[42][7];
              muxOutConnector[35] = fifoOut[43][7];
              muxOutConnector[36] = fifoOut[44][7];
              muxOutConnector[37] = fifoOut[45][7];
              muxOutConnector[38] = fifoOut[46][7];
              muxOutConnector[39] = fifoOut[47][7];
              muxOutConnector[40] = fifoOut[48][7];
              muxOutConnector[41] = fifoOut[49][7];
              muxOutConnector[42] = fifoOut[50][7];
              muxOutConnector[43] = fifoOut[51][7];
              muxOutConnector[44] = fifoOut[26][6];
              muxOutConnector[45] = fifoOut[27][6];
              muxOutConnector[46] = fifoOut[28][6];
              muxOutConnector[47] = fifoOut[29][6];
              muxOutConnector[48] = fifoOut[30][6];
              muxOutConnector[49] = fifoOut[31][6];
              muxOutConnector[50] = fifoOut[32][6];
              muxOutConnector[51] = fifoOut[33][6];
         end
         13: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[43][15];
              muxOutConnector[9] = fifoOut[44][15];
              muxOutConnector[10] = fifoOut[45][15];
              muxOutConnector[11] = fifoOut[46][15];
              muxOutConnector[12] = fifoOut[47][15];
              muxOutConnector[13] = fifoOut[48][15];
              muxOutConnector[14] = fifoOut[49][15];
              muxOutConnector[15] = fifoOut[50][15];
              muxOutConnector[16] = fifoOut[51][15];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][7];
              muxOutConnector[27] = fifoOut[35][7];
              muxOutConnector[28] = fifoOut[36][7];
              muxOutConnector[29] = fifoOut[37][7];
              muxOutConnector[30] = fifoOut[38][7];
              muxOutConnector[31] = fifoOut[39][7];
              muxOutConnector[32] = fifoOut[40][7];
              muxOutConnector[33] = fifoOut[41][7];
              muxOutConnector[34] = fifoOut[42][7];
              muxOutConnector[35] = fifoOut[43][7];
              muxOutConnector[36] = fifoOut[44][7];
              muxOutConnector[37] = fifoOut[45][7];
              muxOutConnector[38] = fifoOut[46][7];
              muxOutConnector[39] = fifoOut[47][7];
              muxOutConnector[40] = fifoOut[48][7];
              muxOutConnector[41] = fifoOut[49][7];
              muxOutConnector[42] = fifoOut[50][7];
              muxOutConnector[43] = fifoOut[51][7];
              muxOutConnector[44] = fifoOut[26][6];
              muxOutConnector[45] = fifoOut[27][6];
              muxOutConnector[46] = fifoOut[28][6];
              muxOutConnector[47] = fifoOut[29][6];
              muxOutConnector[48] = fifoOut[30][6];
              muxOutConnector[49] = fifoOut[31][6];
              muxOutConnector[50] = fifoOut[32][6];
              muxOutConnector[51] = fifoOut[33][6];
         end
         14: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[43][15];
              muxOutConnector[9] = fifoOut[44][15];
              muxOutConnector[10] = fifoOut[45][15];
              muxOutConnector[11] = fifoOut[46][15];
              muxOutConnector[12] = fifoOut[47][15];
              muxOutConnector[13] = fifoOut[48][15];
              muxOutConnector[14] = fifoOut[49][15];
              muxOutConnector[15] = fifoOut[50][15];
              muxOutConnector[16] = fifoOut[51][15];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][7];
              muxOutConnector[27] = fifoOut[35][7];
              muxOutConnector[28] = fifoOut[36][7];
              muxOutConnector[29] = fifoOut[37][7];
              muxOutConnector[30] = fifoOut[38][7];
              muxOutConnector[31] = fifoOut[39][7];
              muxOutConnector[32] = fifoOut[40][7];
              muxOutConnector[33] = fifoOut[41][7];
              muxOutConnector[34] = fifoOut[42][7];
              muxOutConnector[35] = fifoOut[43][7];
              muxOutConnector[36] = fifoOut[44][7];
              muxOutConnector[37] = fifoOut[45][7];
              muxOutConnector[38] = fifoOut[46][7];
              muxOutConnector[39] = fifoOut[47][7];
              muxOutConnector[40] = fifoOut[48][7];
              muxOutConnector[41] = fifoOut[49][7];
              muxOutConnector[42] = fifoOut[50][7];
              muxOutConnector[43] = fifoOut[51][7];
              muxOutConnector[44] = fifoOut[26][6];
              muxOutConnector[45] = fifoOut[27][6];
              muxOutConnector[46] = fifoOut[28][6];
              muxOutConnector[47] = fifoOut[29][6];
              muxOutConnector[48] = fifoOut[30][6];
              muxOutConnector[49] = fifoOut[31][6];
              muxOutConnector[50] = fifoOut[32][6];
              muxOutConnector[51] = fifoOut[33][6];
         end
         15: begin
              muxOutConnector[0] = fifoOut[35][15];
              muxOutConnector[1] = fifoOut[36][15];
              muxOutConnector[2] = fifoOut[37][15];
              muxOutConnector[3] = fifoOut[38][15];
              muxOutConnector[4] = fifoOut[39][15];
              muxOutConnector[5] = fifoOut[40][15];
              muxOutConnector[6] = fifoOut[41][15];
              muxOutConnector[7] = fifoOut[42][15];
              muxOutConnector[8] = fifoOut[19][12];
              muxOutConnector[9] = fifoOut[20][12];
              muxOutConnector[10] = fifoOut[21][12];
              muxOutConnector[11] = fifoOut[22][12];
              muxOutConnector[12] = fifoOut[23][12];
              muxOutConnector[13] = fifoOut[24][12];
              muxOutConnector[14] = fifoOut[25][12];
              muxOutConnector[15] = fifoOut[0][11];
              muxOutConnector[16] = fifoOut[1][11];
              muxOutConnector[17] = fifoOut[2][11];
              muxOutConnector[18] = fifoOut[3][11];
              muxOutConnector[19] = fifoOut[4][11];
              muxOutConnector[20] = fifoOut[5][11];
              muxOutConnector[21] = fifoOut[6][11];
              muxOutConnector[22] = fifoOut[7][11];
              muxOutConnector[23] = fifoOut[8][11];
              muxOutConnector[24] = fifoOut[9][11];
              muxOutConnector[25] = fifoOut[10][11];
              muxOutConnector[26] = fifoOut[34][7];
              muxOutConnector[27] = fifoOut[35][7];
              muxOutConnector[28] = fifoOut[36][7];
              muxOutConnector[29] = fifoOut[37][7];
              muxOutConnector[30] = fifoOut[38][7];
              muxOutConnector[31] = fifoOut[39][7];
              muxOutConnector[32] = fifoOut[40][7];
              muxOutConnector[33] = fifoOut[41][7];
              muxOutConnector[34] = fifoOut[42][7];
              muxOutConnector[35] = fifoOut[43][7];
              muxOutConnector[36] = fifoOut[44][7];
              muxOutConnector[37] = fifoOut[45][7];
              muxOutConnector[38] = fifoOut[46][7];
              muxOutConnector[39] = fifoOut[47][7];
              muxOutConnector[40] = fifoOut[48][7];
              muxOutConnector[41] = fifoOut[49][7];
              muxOutConnector[42] = fifoOut[50][7];
              muxOutConnector[43] = fifoOut[51][7];
              muxOutConnector[44] = fifoOut[26][6];
              muxOutConnector[45] = fifoOut[27][6];
              muxOutConnector[46] = fifoOut[28][6];
              muxOutConnector[47] = fifoOut[29][6];
              muxOutConnector[48] = fifoOut[30][6];
              muxOutConnector[49] = fifoOut[31][6];
              muxOutConnector[50] = fifoOut[32][6];
              muxOutConnector[51] = fifoOut[33][6];
         end
         16: begin
              muxOutConnector[0] = fifoOut[11][12];
              muxOutConnector[1] = fifoOut[12][12];
              muxOutConnector[2] = fifoOut[13][12];
              muxOutConnector[3] = fifoOut[14][12];
              muxOutConnector[4] = fifoOut[15][12];
              muxOutConnector[5] = fifoOut[16][12];
              muxOutConnector[6] = fifoOut[17][12];
              muxOutConnector[7] = fifoOut[18][12];
              muxOutConnector[8] = fifoOut[19][12];
              muxOutConnector[9] = fifoOut[20][12];
              muxOutConnector[10] = fifoOut[21][12];
              muxOutConnector[11] = fifoOut[22][12];
              muxOutConnector[12] = fifoOut[23][12];
              muxOutConnector[13] = fifoOut[24][12];
              muxOutConnector[14] = fifoOut[25][12];
              muxOutConnector[15] = fifoOut[0][11];
              muxOutConnector[16] = fifoOut[1][11];
              muxOutConnector[17] = fifoOut[2][11];
              muxOutConnector[18] = fifoOut[3][11];
              muxOutConnector[19] = fifoOut[4][11];
              muxOutConnector[20] = fifoOut[5][11];
              muxOutConnector[21] = fifoOut[6][11];
              muxOutConnector[22] = fifoOut[7][11];
              muxOutConnector[23] = fifoOut[8][11];
              muxOutConnector[24] = fifoOut[9][11];
              muxOutConnector[25] = fifoOut[10][11];
              muxOutConnector[26] = fifoOut[34][7];
              muxOutConnector[27] = fifoOut[35][7];
              muxOutConnector[28] = fifoOut[36][7];
              muxOutConnector[29] = fifoOut[37][7];
              muxOutConnector[30] = fifoOut[38][7];
              muxOutConnector[31] = fifoOut[39][7];
              muxOutConnector[32] = fifoOut[40][7];
              muxOutConnector[33] = fifoOut[41][7];
              muxOutConnector[34] = fifoOut[42][7];
              muxOutConnector[35] = fifoOut[43][7];
              muxOutConnector[36] = fifoOut[44][7];
              muxOutConnector[37] = fifoOut[45][7];
              muxOutConnector[38] = fifoOut[46][7];
              muxOutConnector[39] = fifoOut[47][7];
              muxOutConnector[40] = fifoOut[48][7];
              muxOutConnector[41] = fifoOut[49][7];
              muxOutConnector[42] = fifoOut[50][7];
              muxOutConnector[43] = fifoOut[51][7];
              muxOutConnector[44] = fifoOut[26][6];
              muxOutConnector[45] = fifoOut[27][6];
              muxOutConnector[46] = fifoOut[28][6];
              muxOutConnector[47] = fifoOut[29][6];
              muxOutConnector[48] = fifoOut[30][6];
              muxOutConnector[49] = fifoOut[31][6];
              muxOutConnector[50] = fifoOut[32][6];
              muxOutConnector[51] = fifoOut[33][6];
         end
         17: begin
              muxOutConnector[0] = fifoOut[11][12];
              muxOutConnector[1] = fifoOut[12][12];
              muxOutConnector[2] = fifoOut[13][12];
              muxOutConnector[3] = fifoOut[14][12];
              muxOutConnector[4] = fifoOut[15][12];
              muxOutConnector[5] = fifoOut[16][12];
              muxOutConnector[6] = fifoOut[17][12];
              muxOutConnector[7] = fifoOut[18][12];
              muxOutConnector[8] = fifoOut[19][12];
              muxOutConnector[9] = fifoOut[20][12];
              muxOutConnector[10] = fifoOut[21][12];
              muxOutConnector[11] = fifoOut[22][12];
              muxOutConnector[12] = fifoOut[23][12];
              muxOutConnector[13] = fifoOut[24][12];
              muxOutConnector[14] = fifoOut[25][12];
              muxOutConnector[15] = fifoOut[0][11];
              muxOutConnector[16] = fifoOut[1][11];
              muxOutConnector[17] = fifoOut[2][11];
              muxOutConnector[18] = fifoOut[3][11];
              muxOutConnector[19] = fifoOut[4][11];
              muxOutConnector[20] = fifoOut[5][11];
              muxOutConnector[21] = fifoOut[6][11];
              muxOutConnector[22] = fifoOut[7][11];
              muxOutConnector[23] = fifoOut[8][11];
              muxOutConnector[24] = fifoOut[9][11];
              muxOutConnector[25] = fifoOut[10][11];
              muxOutConnector[26] = fifoOut[34][7];
              muxOutConnector[27] = fifoOut[35][7];
              muxOutConnector[28] = fifoOut[36][7];
              muxOutConnector[29] = fifoOut[37][7];
              muxOutConnector[30] = fifoOut[38][7];
              muxOutConnector[31] = fifoOut[39][7];
              muxOutConnector[32] = fifoOut[40][7];
              muxOutConnector[33] = fifoOut[41][7];
              muxOutConnector[34] = fifoOut[42][7];
              muxOutConnector[35] = fifoOut[43][7];
              muxOutConnector[36] = fifoOut[44][7];
              muxOutConnector[37] = fifoOut[45][7];
              muxOutConnector[38] = fifoOut[46][7];
              muxOutConnector[39] = fifoOut[47][7];
              muxOutConnector[40] = fifoOut[48][7];
              muxOutConnector[41] = fifoOut[49][7];
              muxOutConnector[42] = fifoOut[50][7];
              muxOutConnector[43] = fifoOut[51][7];
              muxOutConnector[44] = fifoOut[26][6];
              muxOutConnector[45] = fifoOut[27][6];
              muxOutConnector[46] = fifoOut[28][6];
              muxOutConnector[47] = fifoOut[29][6];
              muxOutConnector[48] = fifoOut[30][6];
              muxOutConnector[49] = fifoOut[31][6];
              muxOutConnector[50] = fifoOut[32][6];
              muxOutConnector[51] = fifoOut[33][6];
         end
         18: begin
              muxOutConnector[0] = fifoOut[11][12];
              muxOutConnector[1] = fifoOut[12][12];
              muxOutConnector[2] = fifoOut[13][12];
              muxOutConnector[3] = fifoOut[14][12];
              muxOutConnector[4] = fifoOut[15][12];
              muxOutConnector[5] = fifoOut[16][12];
              muxOutConnector[6] = fifoOut[17][12];
              muxOutConnector[7] = fifoOut[18][12];
              muxOutConnector[8] = fifoOut[19][12];
              muxOutConnector[9] = fifoOut[20][12];
              muxOutConnector[10] = fifoOut[21][12];
              muxOutConnector[11] = fifoOut[22][12];
              muxOutConnector[12] = fifoOut[23][12];
              muxOutConnector[13] = fifoOut[24][12];
              muxOutConnector[14] = fifoOut[25][12];
              muxOutConnector[15] = fifoOut[0][11];
              muxOutConnector[16] = fifoOut[1][11];
              muxOutConnector[17] = fifoOut[2][11];
              muxOutConnector[18] = fifoOut[3][11];
              muxOutConnector[19] = fifoOut[4][11];
              muxOutConnector[20] = fifoOut[5][11];
              muxOutConnector[21] = fifoOut[6][11];
              muxOutConnector[22] = fifoOut[7][11];
              muxOutConnector[23] = fifoOut[8][11];
              muxOutConnector[24] = fifoOut[9][11];
              muxOutConnector[25] = fifoOut[10][11];
              muxOutConnector[26] = fifoOut[34][7];
              muxOutConnector[27] = fifoOut[35][7];
              muxOutConnector[28] = fifoOut[36][7];
              muxOutConnector[29] = fifoOut[37][7];
              muxOutConnector[30] = fifoOut[38][7];
              muxOutConnector[31] = fifoOut[39][7];
              muxOutConnector[32] = fifoOut[40][7];
              muxOutConnector[33] = fifoOut[41][7];
              muxOutConnector[34] = fifoOut[42][7];
              muxOutConnector[35] = fifoOut[43][7];
              muxOutConnector[36] = fifoOut[44][7];
              muxOutConnector[37] = fifoOut[45][7];
              muxOutConnector[38] = fifoOut[46][7];
              muxOutConnector[39] = fifoOut[47][7];
              muxOutConnector[40] = fifoOut[48][7];
              muxOutConnector[41] = fifoOut[49][7];
              muxOutConnector[42] = fifoOut[50][7];
              muxOutConnector[43] = fifoOut[51][7];
              muxOutConnector[44] = fifoOut[26][6];
              muxOutConnector[45] = fifoOut[27][6];
              muxOutConnector[46] = fifoOut[28][6];
              muxOutConnector[47] = fifoOut[29][6];
              muxOutConnector[48] = fifoOut[30][6];
              muxOutConnector[49] = fifoOut[31][6];
              muxOutConnector[50] = fifoOut[32][6];
              muxOutConnector[51] = fifoOut[33][6];
         end
         19: begin
              muxOutConnector[0] = fifoOut[11][12];
              muxOutConnector[1] = fifoOut[12][12];
              muxOutConnector[2] = fifoOut[13][12];
              muxOutConnector[3] = fifoOut[14][12];
              muxOutConnector[4] = fifoOut[15][12];
              muxOutConnector[5] = fifoOut[16][12];
              muxOutConnector[6] = fifoOut[17][12];
              muxOutConnector[7] = fifoOut[18][12];
              muxOutConnector[8] = fifoOut[19][12];
              muxOutConnector[9] = fifoOut[20][12];
              muxOutConnector[10] = fifoOut[21][12];
              muxOutConnector[11] = fifoOut[22][12];
              muxOutConnector[12] = fifoOut[23][12];
              muxOutConnector[13] = fifoOut[24][12];
              muxOutConnector[14] = fifoOut[25][12];
              muxOutConnector[15] = fifoOut[0][11];
              muxOutConnector[16] = fifoOut[1][11];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[34][7];
              muxOutConnector[27] = fifoOut[35][7];
              muxOutConnector[28] = fifoOut[36][7];
              muxOutConnector[29] = fifoOut[37][7];
              muxOutConnector[30] = fifoOut[38][7];
              muxOutConnector[31] = fifoOut[39][7];
              muxOutConnector[32] = fifoOut[40][7];
              muxOutConnector[33] = fifoOut[41][7];
              muxOutConnector[34] = fifoOut[42][7];
              muxOutConnector[35] = fifoOut[43][7];
              muxOutConnector[36] = fifoOut[44][7];
              muxOutConnector[37] = fifoOut[45][7];
              muxOutConnector[38] = fifoOut[46][7];
              muxOutConnector[39] = fifoOut[47][7];
              muxOutConnector[40] = fifoOut[48][7];
              muxOutConnector[41] = fifoOut[49][7];
              muxOutConnector[42] = fifoOut[50][7];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
         end
         default: begin
               for(i=0;i<muxOutSymbols;i=i+1)begin
                muxOutConnector[i] = 0;
              end
         end
//hgjhgbuiguigbigbgbgbui
         endcase
    end
endcase
             end
        endmodule