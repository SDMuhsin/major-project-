`timescale 1ns / 1ps
module LMem0To1_511_circ10_ys_scripted(
        muxOut,
        ly0In,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 13;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            fifoOut[i][0] <= ly0InConnector[i];
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[36][4];
              muxOutConnector[1] = fifoOut[37][4];
              muxOutConnector[2] = fifoOut[38][4];
              muxOutConnector[3] = fifoOut[39][4];
              muxOutConnector[4] = fifoOut[40][4];
              muxOutConnector[5] = fifoOut[41][4];
              muxOutConnector[6] = fifoOut[42][4];
              muxOutConnector[7] = fifoOut[43][4];
              muxOutConnector[8] = fifoOut[44][4];
              muxOutConnector[9] = fifoOut[45][4];
              muxOutConnector[10] = fifoOut[46][4];
              muxOutConnector[11] = fifoOut[47][4];
              muxOutConnector[12] = fifoOut[48][4];
              muxOutConnector[13] = fifoOut[49][4];
              muxOutConnector[14] = fifoOut[50][4];
              muxOutConnector[15] = fifoOut[51][4];
              muxOutConnector[16] = fifoOut[26][3];
              muxOutConnector[17] = fifoOut[27][3];
              muxOutConnector[18] = fifoOut[28][3];
              muxOutConnector[19] = fifoOut[29][3];
              muxOutConnector[20] = fifoOut[30][3];
              muxOutConnector[21] = fifoOut[31][3];
              muxOutConnector[22] = fifoOut[32][3];
              muxOutConnector[23] = fifoOut[33][3];
              muxOutConnector[24] = fifoOut[34][3];
              muxOutConnector[25] = fifoOut[35][3];
              muxOutConnector[26] = fifoOut[15][5];
              muxOutConnector[27] = fifoOut[16][5];
              muxOutConnector[28] = fifoOut[17][5];
              muxOutConnector[29] = fifoOut[18][5];
              muxOutConnector[30] = fifoOut[19][5];
              muxOutConnector[31] = fifoOut[20][5];
              muxOutConnector[32] = fifoOut[21][5];
              muxOutConnector[33] = fifoOut[22][5];
              muxOutConnector[34] = fifoOut[23][5];
              muxOutConnector[35] = fifoOut[24][5];
              muxOutConnector[36] = fifoOut[26][12];
              muxOutConnector[37] = fifoOut[27][12];
              muxOutConnector[38] = fifoOut[28][12];
              muxOutConnector[39] = fifoOut[29][12];
              muxOutConnector[40] = fifoOut[30][12];
              muxOutConnector[41] = fifoOut[31][12];
              muxOutConnector[42] = fifoOut[32][12];
              muxOutConnector[43] = fifoOut[33][12];
              muxOutConnector[44] = fifoOut[34][12];
              muxOutConnector[45] = fifoOut[35][12];
              muxOutConnector[46] = fifoOut[36][12];
              muxOutConnector[47] = fifoOut[37][12];
              muxOutConnector[48] = fifoOut[38][12];
              muxOutConnector[49] = fifoOut[39][12];
              muxOutConnector[50] = fifoOut[40][12];
              muxOutConnector[51] = fifoOut[41][12];
       end
       1: begin
              muxOutConnector[0] = fifoOut[36][4];
              muxOutConnector[1] = fifoOut[37][4];
              muxOutConnector[2] = fifoOut[38][4];
              muxOutConnector[3] = fifoOut[39][4];
              muxOutConnector[4] = fifoOut[40][4];
              muxOutConnector[5] = fifoOut[41][4];
              muxOutConnector[6] = fifoOut[42][4];
              muxOutConnector[7] = fifoOut[43][4];
              muxOutConnector[8] = fifoOut[44][4];
              muxOutConnector[9] = fifoOut[45][4];
              muxOutConnector[10] = fifoOut[46][4];
              muxOutConnector[11] = fifoOut[47][4];
              muxOutConnector[12] = fifoOut[48][4];
              muxOutConnector[13] = fifoOut[49][4];
              muxOutConnector[14] = fifoOut[50][4];
              muxOutConnector[15] = fifoOut[51][4];
              muxOutConnector[16] = fifoOut[26][3];
              muxOutConnector[17] = fifoOut[27][3];
              muxOutConnector[18] = fifoOut[28][3];
              muxOutConnector[19] = fifoOut[29][3];
              muxOutConnector[20] = fifoOut[30][3];
              muxOutConnector[21] = fifoOut[31][3];
              muxOutConnector[22] = fifoOut[32][3];
              muxOutConnector[23] = fifoOut[33][3];
              muxOutConnector[24] = fifoOut[34][3];
              muxOutConnector[25] = fifoOut[35][3];
              muxOutConnector[26] = fifoOut[15][5];
              muxOutConnector[27] = fifoOut[16][5];
              muxOutConnector[28] = fifoOut[17][5];
              muxOutConnector[29] = fifoOut[18][5];
              muxOutConnector[30] = fifoOut[19][5];
              muxOutConnector[31] = fifoOut[20][5];
              muxOutConnector[32] = fifoOut[21][5];
              muxOutConnector[33] = fifoOut[22][5];
              muxOutConnector[34] = fifoOut[23][5];
              muxOutConnector[35] = fifoOut[24][5];
              muxOutConnector[36] = fifoOut[26][12];
              muxOutConnector[37] = fifoOut[27][12];
              muxOutConnector[38] = fifoOut[28][12];
              muxOutConnector[39] = fifoOut[29][12];
              muxOutConnector[40] = fifoOut[30][12];
              muxOutConnector[41] = fifoOut[31][12];
              muxOutConnector[42] = fifoOut[32][12];
              muxOutConnector[43] = fifoOut[33][12];
              muxOutConnector[44] = fifoOut[34][12];
              muxOutConnector[45] = fifoOut[35][12];
              muxOutConnector[46] = fifoOut[36][12];
              muxOutConnector[47] = fifoOut[37][12];
              muxOutConnector[48] = fifoOut[38][12];
              muxOutConnector[49] = fifoOut[39][12];
              muxOutConnector[50] = fifoOut[40][12];
              muxOutConnector[51] = fifoOut[41][12];
       end
       2: begin
              muxOutConnector[0] = fifoOut[36][4];
              muxOutConnector[1] = fifoOut[37][4];
              muxOutConnector[2] = fifoOut[38][4];
              muxOutConnector[3] = fifoOut[39][4];
              muxOutConnector[4] = fifoOut[40][4];
              muxOutConnector[5] = fifoOut[41][4];
              muxOutConnector[6] = fifoOut[42][4];
              muxOutConnector[7] = fifoOut[43][4];
              muxOutConnector[8] = fifoOut[44][4];
              muxOutConnector[9] = fifoOut[45][4];
              muxOutConnector[10] = fifoOut[46][4];
              muxOutConnector[11] = fifoOut[47][4];
              muxOutConnector[12] = fifoOut[48][4];
              muxOutConnector[13] = fifoOut[49][4];
              muxOutConnector[14] = fifoOut[50][4];
              muxOutConnector[15] = fifoOut[51][4];
              muxOutConnector[16] = fifoOut[26][3];
              muxOutConnector[17] = fifoOut[27][3];
              muxOutConnector[18] = fifoOut[28][3];
              muxOutConnector[19] = fifoOut[29][3];
              muxOutConnector[20] = fifoOut[30][3];
              muxOutConnector[21] = fifoOut[31][3];
              muxOutConnector[22] = fifoOut[32][3];
              muxOutConnector[23] = fifoOut[33][3];
              muxOutConnector[24] = fifoOut[34][3];
              muxOutConnector[25] = fifoOut[35][3];
              muxOutConnector[26] = fifoOut[15][5];
              muxOutConnector[27] = fifoOut[16][5];
              muxOutConnector[28] = fifoOut[17][5];
              muxOutConnector[29] = fifoOut[18][5];
              muxOutConnector[30] = fifoOut[19][5];
              muxOutConnector[31] = fifoOut[20][5];
              muxOutConnector[32] = fifoOut[21][5];
              muxOutConnector[33] = fifoOut[22][5];
              muxOutConnector[34] = fifoOut[23][5];
              muxOutConnector[35] = fifoOut[24][5];
              muxOutConnector[36] = fifoOut[26][12];
              muxOutConnector[37] = fifoOut[27][12];
              muxOutConnector[38] = fifoOut[28][12];
              muxOutConnector[39] = fifoOut[29][12];
              muxOutConnector[40] = fifoOut[30][12];
              muxOutConnector[41] = fifoOut[31][12];
              muxOutConnector[42] = fifoOut[32][12];
              muxOutConnector[43] = fifoOut[33][12];
              muxOutConnector[44] = fifoOut[34][12];
              muxOutConnector[45] = fifoOut[35][12];
              muxOutConnector[46] = fifoOut[36][12];
              muxOutConnector[47] = fifoOut[37][12];
              muxOutConnector[48] = fifoOut[38][12];
              muxOutConnector[49] = fifoOut[39][12];
              muxOutConnector[50] = fifoOut[40][12];
              muxOutConnector[51] = fifoOut[41][12];
       end
       3: begin
              muxOutConnector[0] = fifoOut[36][4];
              muxOutConnector[1] = fifoOut[37][4];
              muxOutConnector[2] = fifoOut[38][4];
              muxOutConnector[3] = fifoOut[39][4];
              muxOutConnector[4] = fifoOut[40][4];
              muxOutConnector[5] = fifoOut[41][4];
              muxOutConnector[6] = fifoOut[42][4];
              muxOutConnector[7] = fifoOut[43][4];
              muxOutConnector[8] = fifoOut[44][4];
              muxOutConnector[9] = fifoOut[45][4];
              muxOutConnector[10] = fifoOut[46][4];
              muxOutConnector[11] = fifoOut[47][4];
              muxOutConnector[12] = fifoOut[48][4];
              muxOutConnector[13] = fifoOut[49][4];
              muxOutConnector[14] = fifoOut[50][4];
              muxOutConnector[15] = fifoOut[51][4];
              muxOutConnector[16] = fifoOut[26][3];
              muxOutConnector[17] = fifoOut[27][3];
              muxOutConnector[18] = fifoOut[28][3];
              muxOutConnector[19] = fifoOut[29][3];
              muxOutConnector[20] = fifoOut[30][3];
              muxOutConnector[21] = fifoOut[31][3];
              muxOutConnector[22] = fifoOut[32][3];
              muxOutConnector[23] = fifoOut[33][3];
              muxOutConnector[24] = fifoOut[34][3];
              muxOutConnector[25] = fifoOut[35][3];
              muxOutConnector[26] = fifoOut[15][5];
              muxOutConnector[27] = fifoOut[16][5];
              muxOutConnector[28] = fifoOut[17][5];
              muxOutConnector[29] = fifoOut[18][5];
              muxOutConnector[30] = fifoOut[19][5];
              muxOutConnector[31] = fifoOut[20][5];
              muxOutConnector[32] = fifoOut[21][5];
              muxOutConnector[33] = fifoOut[22][5];
              muxOutConnector[34] = fifoOut[23][5];
              muxOutConnector[35] = fifoOut[24][5];
              muxOutConnector[36] = fifoOut[26][12];
              muxOutConnector[37] = fifoOut[27][12];
              muxOutConnector[38] = fifoOut[28][12];
              muxOutConnector[39] = fifoOut[29][12];
              muxOutConnector[40] = fifoOut[30][12];
              muxOutConnector[41] = fifoOut[31][12];
              muxOutConnector[42] = fifoOut[32][12];
              muxOutConnector[43] = fifoOut[33][12];
              muxOutConnector[44] = fifoOut[34][12];
              muxOutConnector[45] = fifoOut[35][12];
              muxOutConnector[46] = fifoOut[36][12];
              muxOutConnector[47] = fifoOut[37][12];
              muxOutConnector[48] = fifoOut[38][12];
              muxOutConnector[49] = fifoOut[39][12];
              muxOutConnector[50] = fifoOut[40][12];
              muxOutConnector[51] = fifoOut[41][12];
       end
       4: begin
              muxOutConnector[0] = fifoOut[36][4];
              muxOutConnector[1] = fifoOut[37][4];
              muxOutConnector[2] = fifoOut[38][4];
              muxOutConnector[3] = fifoOut[39][4];
              muxOutConnector[4] = fifoOut[40][4];
              muxOutConnector[5] = fifoOut[41][4];
              muxOutConnector[6] = fifoOut[42][4];
              muxOutConnector[7] = fifoOut[25][3];
              muxOutConnector[8] = fifoOut[0][2];
              muxOutConnector[9] = fifoOut[1][2];
              muxOutConnector[10] = fifoOut[2][2];
              muxOutConnector[11] = fifoOut[3][2];
              muxOutConnector[12] = fifoOut[4][2];
              muxOutConnector[13] = fifoOut[5][2];
              muxOutConnector[14] = fifoOut[6][2];
              muxOutConnector[15] = fifoOut[7][2];
              muxOutConnector[16] = fifoOut[8][2];
              muxOutConnector[17] = fifoOut[9][2];
              muxOutConnector[18] = fifoOut[10][2];
              muxOutConnector[19] = fifoOut[11][2];
              muxOutConnector[20] = fifoOut[12][2];
              muxOutConnector[21] = fifoOut[13][2];
              muxOutConnector[22] = fifoOut[14][2];
              muxOutConnector[23] = fifoOut[15][2];
              muxOutConnector[24] = fifoOut[16][2];
              muxOutConnector[25] = fifoOut[17][2];
              muxOutConnector[26] = fifoOut[15][5];
              muxOutConnector[27] = fifoOut[16][5];
              muxOutConnector[28] = fifoOut[17][5];
              muxOutConnector[29] = fifoOut[18][5];
              muxOutConnector[30] = fifoOut[19][5];
              muxOutConnector[31] = fifoOut[20][5];
              muxOutConnector[32] = fifoOut[21][5];
              muxOutConnector[33] = fifoOut[22][5];
              muxOutConnector[34] = fifoOut[23][5];
              muxOutConnector[35] = fifoOut[24][5];
              muxOutConnector[36] = fifoOut[26][12];
              muxOutConnector[37] = fifoOut[27][12];
              muxOutConnector[38] = fifoOut[28][12];
              muxOutConnector[39] = fifoOut[29][12];
              muxOutConnector[40] = fifoOut[30][12];
              muxOutConnector[41] = fifoOut[31][12];
              muxOutConnector[42] = fifoOut[32][12];
              muxOutConnector[43] = fifoOut[33][12];
              muxOutConnector[44] = fifoOut[34][12];
              muxOutConnector[45] = fifoOut[35][12];
              muxOutConnector[46] = fifoOut[36][12];
              muxOutConnector[47] = fifoOut[37][12];
              muxOutConnector[48] = fifoOut[38][12];
              muxOutConnector[49] = fifoOut[39][12];
              muxOutConnector[50] = fifoOut[40][12];
              muxOutConnector[51] = fifoOut[41][12];
       end
       5: begin
              muxOutConnector[0] = fifoOut[18][3];
              muxOutConnector[1] = fifoOut[19][3];
              muxOutConnector[2] = fifoOut[20][3];
              muxOutConnector[3] = fifoOut[21][3];
              muxOutConnector[4] = fifoOut[22][3];
              muxOutConnector[5] = fifoOut[23][3];
              muxOutConnector[6] = fifoOut[24][3];
              muxOutConnector[7] = fifoOut[25][3];
              muxOutConnector[8] = fifoOut[0][2];
              muxOutConnector[9] = fifoOut[1][2];
              muxOutConnector[10] = fifoOut[2][2];
              muxOutConnector[11] = fifoOut[3][2];
              muxOutConnector[12] = fifoOut[4][2];
              muxOutConnector[13] = fifoOut[5][2];
              muxOutConnector[14] = fifoOut[6][2];
              muxOutConnector[15] = fifoOut[7][2];
              muxOutConnector[16] = fifoOut[8][2];
              muxOutConnector[17] = fifoOut[9][2];
              muxOutConnector[18] = fifoOut[10][2];
              muxOutConnector[19] = fifoOut[11][2];
              muxOutConnector[20] = fifoOut[12][2];
              muxOutConnector[21] = fifoOut[13][2];
              muxOutConnector[22] = fifoOut[14][2];
              muxOutConnector[23] = fifoOut[15][2];
              muxOutConnector[24] = fifoOut[16][2];
              muxOutConnector[25] = fifoOut[17][2];
              muxOutConnector[26] = fifoOut[15][5];
              muxOutConnector[27] = fifoOut[16][5];
              muxOutConnector[28] = fifoOut[44][0];
              muxOutConnector[29] = fifoOut[45][0];
              muxOutConnector[30] = fifoOut[46][0];
              muxOutConnector[31] = fifoOut[47][0];
              muxOutConnector[32] = fifoOut[48][0];
              muxOutConnector[33] = fifoOut[49][0];
              muxOutConnector[34] = fifoOut[50][0];
              muxOutConnector[35] = fifoOut[51][0];
              muxOutConnector[36] = fifoOut[26][12];
              muxOutConnector[37] = fifoOut[27][12];
              muxOutConnector[38] = fifoOut[28][12];
              muxOutConnector[39] = fifoOut[29][12];
              muxOutConnector[40] = fifoOut[30][12];
              muxOutConnector[41] = fifoOut[31][12];
              muxOutConnector[42] = fifoOut[32][12];
              muxOutConnector[43] = fifoOut[33][12];
              muxOutConnector[44] = fifoOut[34][12];
              muxOutConnector[45] = fifoOut[35][12];
              muxOutConnector[46] = fifoOut[36][12];
              muxOutConnector[47] = fifoOut[37][12];
              muxOutConnector[48] = fifoOut[38][12];
              muxOutConnector[49] = fifoOut[39][12];
              muxOutConnector[50] = fifoOut[40][12];
              muxOutConnector[51] = fifoOut[41][12];
       end
       6: begin
              muxOutConnector[0] = fifoOut[18][3];
              muxOutConnector[1] = fifoOut[19][3];
              muxOutConnector[2] = fifoOut[20][3];
              muxOutConnector[3] = fifoOut[21][3];
              muxOutConnector[4] = fifoOut[22][3];
              muxOutConnector[5] = fifoOut[23][3];
              muxOutConnector[6] = fifoOut[24][3];
              muxOutConnector[7] = fifoOut[25][3];
              muxOutConnector[8] = fifoOut[0][2];
              muxOutConnector[9] = fifoOut[1][2];
              muxOutConnector[10] = fifoOut[2][2];
              muxOutConnector[11] = fifoOut[3][2];
              muxOutConnector[12] = fifoOut[4][2];
              muxOutConnector[13] = fifoOut[5][2];
              muxOutConnector[14] = fifoOut[6][2];
              muxOutConnector[15] = fifoOut[7][2];
              muxOutConnector[16] = fifoOut[8][2];
              muxOutConnector[17] = fifoOut[9][2];
              muxOutConnector[18] = fifoOut[10][2];
              muxOutConnector[19] = fifoOut[11][2];
              muxOutConnector[20] = fifoOut[12][2];
              muxOutConnector[21] = fifoOut[13][2];
              muxOutConnector[22] = fifoOut[14][2];
              muxOutConnector[23] = fifoOut[15][2];
              muxOutConnector[24] = fifoOut[16][2];
              muxOutConnector[25] = fifoOut[17][2];
              muxOutConnector[26] = fifoOut[42][0];
              muxOutConnector[27] = fifoOut[43][0];
              muxOutConnector[28] = fifoOut[44][0];
              muxOutConnector[29] = fifoOut[45][0];
              muxOutConnector[30] = fifoOut[46][0];
              muxOutConnector[31] = fifoOut[47][0];
              muxOutConnector[32] = fifoOut[48][0];
              muxOutConnector[33] = fifoOut[49][0];
              muxOutConnector[34] = fifoOut[50][0];
              muxOutConnector[35] = fifoOut[51][0];
              muxOutConnector[36] = fifoOut[26][12];
              muxOutConnector[37] = fifoOut[27][12];
              muxOutConnector[38] = fifoOut[28][12];
              muxOutConnector[39] = fifoOut[29][12];
              muxOutConnector[40] = fifoOut[30][12];
              muxOutConnector[41] = fifoOut[31][12];
              muxOutConnector[42] = fifoOut[32][12];
              muxOutConnector[43] = fifoOut[33][12];
              muxOutConnector[44] = fifoOut[34][12];
              muxOutConnector[45] = fifoOut[35][12];
              muxOutConnector[46] = fifoOut[36][12];
              muxOutConnector[47] = fifoOut[37][12];
              muxOutConnector[48] = fifoOut[38][12];
              muxOutConnector[49] = fifoOut[39][12];
              muxOutConnector[50] = fifoOut[40][12];
              muxOutConnector[51] = fifoOut[41][12];
       end
       7: begin
              muxOutConnector[0] = fifoOut[18][3];
              muxOutConnector[1] = fifoOut[19][3];
              muxOutConnector[2] = fifoOut[20][3];
              muxOutConnector[3] = fifoOut[21][3];
              muxOutConnector[4] = fifoOut[22][3];
              muxOutConnector[5] = fifoOut[23][3];
              muxOutConnector[6] = fifoOut[24][3];
              muxOutConnector[7] = fifoOut[25][3];
              muxOutConnector[8] = fifoOut[0][2];
              muxOutConnector[9] = fifoOut[1][2];
              muxOutConnector[10] = fifoOut[2][2];
              muxOutConnector[11] = fifoOut[3][2];
              muxOutConnector[12] = fifoOut[4][2];
              muxOutConnector[13] = fifoOut[5][2];
              muxOutConnector[14] = fifoOut[6][2];
              muxOutConnector[15] = fifoOut[7][2];
              muxOutConnector[16] = fifoOut[8][2];
              muxOutConnector[17] = fifoOut[9][2];
              muxOutConnector[18] = fifoOut[10][2];
              muxOutConnector[19] = fifoOut[11][2];
              muxOutConnector[20] = fifoOut[12][2];
              muxOutConnector[21] = fifoOut[13][2];
              muxOutConnector[22] = fifoOut[14][2];
              muxOutConnector[23] = fifoOut[15][2];
              muxOutConnector[24] = fifoOut[16][2];
              muxOutConnector[25] = fifoOut[17][2];
              muxOutConnector[26] = fifoOut[42][0];
              muxOutConnector[27] = fifoOut[43][0];
              muxOutConnector[28] = fifoOut[44][0];
              muxOutConnector[29] = fifoOut[45][0];
              muxOutConnector[30] = fifoOut[46][0];
              muxOutConnector[31] = fifoOut[47][0];
              muxOutConnector[32] = fifoOut[48][0];
              muxOutConnector[33] = fifoOut[49][0];
              muxOutConnector[34] = fifoOut[50][0];
              muxOutConnector[35] = fifoOut[51][0];
              muxOutConnector[36] = fifoOut[26][12];
              muxOutConnector[37] = fifoOut[27][12];
              muxOutConnector[38] = fifoOut[28][12];
              muxOutConnector[39] = fifoOut[29][12];
              muxOutConnector[40] = fifoOut[30][12];
              muxOutConnector[41] = fifoOut[31][12];
              muxOutConnector[42] = fifoOut[32][12];
              muxOutConnector[43] = fifoOut[33][12];
              muxOutConnector[44] = fifoOut[34][12];
              muxOutConnector[45] = fifoOut[35][12];
              muxOutConnector[46] = fifoOut[36][12];
              muxOutConnector[47] = fifoOut[37][12];
              muxOutConnector[48] = fifoOut[38][12];
              muxOutConnector[49] = fifoOut[39][12];
              muxOutConnector[50] = fifoOut[40][12];
              muxOutConnector[51] = fifoOut[41][12];
       end
       8: begin
              muxOutConnector[0] = fifoOut[18][3];
              muxOutConnector[1] = fifoOut[19][3];
              muxOutConnector[2] = fifoOut[20][3];
              muxOutConnector[3] = fifoOut[21][3];
              muxOutConnector[4] = fifoOut[22][3];
              muxOutConnector[5] = fifoOut[23][3];
              muxOutConnector[6] = fifoOut[24][3];
              muxOutConnector[7] = fifoOut[25][3];
              muxOutConnector[8] = fifoOut[0][2];
              muxOutConnector[9] = fifoOut[1][2];
              muxOutConnector[10] = fifoOut[2][2];
              muxOutConnector[11] = fifoOut[3][2];
              muxOutConnector[12] = fifoOut[4][2];
              muxOutConnector[13] = fifoOut[5][2];
              muxOutConnector[14] = fifoOut[6][2];
              muxOutConnector[15] = fifoOut[7][2];
              muxOutConnector[16] = fifoOut[8][2];
              muxOutConnector[17] = fifoOut[9][2];
              muxOutConnector[18] = fifoOut[10][2];
              muxOutConnector[19] = fifoOut[11][2];
              muxOutConnector[20] = fifoOut[12][2];
              muxOutConnector[21] = fifoOut[13][2];
              muxOutConnector[22] = fifoOut[14][2];
              muxOutConnector[23] = fifoOut[15][2];
              muxOutConnector[24] = fifoOut[16][2];
              muxOutConnector[25] = fifoOut[17][2];
              muxOutConnector[26] = fifoOut[42][0];
              muxOutConnector[27] = fifoOut[43][0];
              muxOutConnector[28] = fifoOut[44][0];
              muxOutConnector[29] = fifoOut[45][0];
              muxOutConnector[30] = fifoOut[46][0];
              muxOutConnector[31] = fifoOut[47][0];
              muxOutConnector[32] = fifoOut[48][0];
              muxOutConnector[33] = fifoOut[49][0];
              muxOutConnector[34] = fifoOut[50][0];
              muxOutConnector[35] = fifoOut[51][0];
              muxOutConnector[36] = fifoOut[26][12];
              muxOutConnector[37] = fifoOut[27][12];
              muxOutConnector[38] = fifoOut[28][12];
              muxOutConnector[39] = fifoOut[29][12];
              muxOutConnector[40] = fifoOut[30][12];
              muxOutConnector[41] = fifoOut[31][12];
              muxOutConnector[42] = fifoOut[32][12];
              muxOutConnector[43] = fifoOut[33][12];
              muxOutConnector[44] = fifoOut[34][12];
              muxOutConnector[45] = fifoOut[35][12];
              muxOutConnector[46] = fifoOut[36][12];
              muxOutConnector[47] = fifoOut[37][12];
              muxOutConnector[48] = fifoOut[38][12];
              muxOutConnector[49] = fifoOut[39][12];
              muxOutConnector[50] = fifoOut[40][12];
              muxOutConnector[51] = fifoOut[41][12];
       end
       9: begin
              muxOutConnector[0] = fifoOut[18][3];
              muxOutConnector[1] = fifoOut[19][3];
              muxOutConnector[2] = fifoOut[20][3];
              muxOutConnector[3] = fifoOut[21][3];
              muxOutConnector[4] = fifoOut[22][3];
              muxOutConnector[5] = fifoOut[23][3];
              muxOutConnector[6] = fifoOut[24][3];
              muxOutConnector[7] = fifoOut[25][3];
              muxOutConnector[8] = fifoOut[0][2];
              muxOutConnector[9] = fifoOut[1][2];
              muxOutConnector[10] = fifoOut[2][2];
              muxOutConnector[11] = fifoOut[3][2];
              muxOutConnector[12] = fifoOut[4][2];
              muxOutConnector[13] = fifoOut[5][2];
              muxOutConnector[14] = fifoOut[6][2];
              muxOutConnector[15] = fifoOut[7][2];
              muxOutConnector[16] = fifoOut[8][2];
              muxOutConnector[17] = fifoOut[9][2];
              muxOutConnector[18] = fifoOut[10][2];
              muxOutConnector[19] = fifoOut[11][2];
              muxOutConnector[20] = fifoOut[12][2];
              muxOutConnector[21] = fifoOut[13][2];
              muxOutConnector[22] = fifoOut[14][2];
              muxOutConnector[23] = fifoOut[15][2];
              muxOutConnector[24] = fifoOut[16][2];
              muxOutConnector[25] = fifoOut[17][2];
              muxOutConnector[26] = fifoOut[42][0];
              muxOutConnector[27] = fifoOut[43][0];
              muxOutConnector[28] = fifoOut[44][0];
              muxOutConnector[29] = fifoOut[45][0];
              muxOutConnector[30] = fifoOut[46][0];
              muxOutConnector[31] = fifoOut[47][0];
              muxOutConnector[32] = fifoOut[48][0];
              muxOutConnector[33] = fifoOut[49][0];
              muxOutConnector[34] = fifoOut[50][0];
              muxOutConnector[35] = fifoOut[51][0];
              muxOutConnector[36] = fifoOut[26][12];
              muxOutConnector[37] = fifoOut[27][12];
              muxOutConnector[38] = fifoOut[28][12];
              muxOutConnector[39] = fifoOut[29][12];
              muxOutConnector[40] = fifoOut[30][12];
              muxOutConnector[41] = fifoOut[31][12];
              muxOutConnector[42] = fifoOut[32][12];
              muxOutConnector[43] = fifoOut[33][12];
              muxOutConnector[44] = fifoOut[34][12];
              muxOutConnector[45] = fifoOut[35][12];
              muxOutConnector[46] = fifoOut[36][12];
              muxOutConnector[47] = fifoOut[37][12];
              muxOutConnector[48] = fifoOut[38][12];
              muxOutConnector[49] = fifoOut[39][12];
              muxOutConnector[50] = fifoOut[40][12];
              muxOutConnector[51] = fifoOut[41][12];
       end
       10: begin
              muxOutConnector[0] = fifoOut[18][3];
              muxOutConnector[1] = fifoOut[19][3];
              muxOutConnector[2] = fifoOut[20][3];
              muxOutConnector[3] = fifoOut[21][3];
              muxOutConnector[4] = fifoOut[22][3];
              muxOutConnector[5] = fifoOut[23][3];
              muxOutConnector[6] = fifoOut[24][3];
              muxOutConnector[7] = fifoOut[25][3];
              muxOutConnector[8] = fifoOut[0][2];
              muxOutConnector[9] = fifoOut[1][2];
              muxOutConnector[10] = fifoOut[2][2];
              muxOutConnector[11] = fifoOut[3][2];
              muxOutConnector[12] = fifoOut[4][2];
              muxOutConnector[13] = fifoOut[5][2];
              muxOutConnector[14] = fifoOut[6][2];
              muxOutConnector[15] = fifoOut[7][2];
              muxOutConnector[16] = fifoOut[8][2];
              muxOutConnector[17] = fifoOut[9][2];
              muxOutConnector[18] = fifoOut[10][2];
              muxOutConnector[19] = fifoOut[11][2];
              muxOutConnector[20] = fifoOut[12][2];
              muxOutConnector[21] = fifoOut[13][2];
              muxOutConnector[22] = fifoOut[14][2];
              muxOutConnector[23] = fifoOut[15][2];
              muxOutConnector[24] = fifoOut[16][2];
              muxOutConnector[25] = fifoOut[17][2];
              muxOutConnector[26] = fifoOut[42][0];
              muxOutConnector[27] = fifoOut[43][0];
              muxOutConnector[28] = fifoOut[44][0];
              muxOutConnector[29] = fifoOut[45][0];
              muxOutConnector[30] = fifoOut[46][0];
              muxOutConnector[31] = fifoOut[47][0];
              muxOutConnector[32] = fifoOut[48][0];
              muxOutConnector[33] = fifoOut[49][0];
              muxOutConnector[34] = fifoOut[50][0];
              muxOutConnector[35] = fifoOut[51][0];
              muxOutConnector[36] = fifoOut[26][12];
              muxOutConnector[37] = fifoOut[27][12];
              muxOutConnector[38] = fifoOut[28][12];
              muxOutConnector[39] = fifoOut[29][12];
              muxOutConnector[40] = fifoOut[30][12];
              muxOutConnector[41] = fifoOut[31][12];
              muxOutConnector[42] = fifoOut[32][12];
              muxOutConnector[43] = fifoOut[33][12];
              muxOutConnector[44] = fifoOut[34][12];
              muxOutConnector[45] = fifoOut[35][12];
              muxOutConnector[46] = fifoOut[36][12];
              muxOutConnector[47] = fifoOut[37][12];
              muxOutConnector[48] = fifoOut[38][12];
              muxOutConnector[49] = fifoOut[39][12];
              muxOutConnector[50] = fifoOut[40][12];
              muxOutConnector[51] = fifoOut[41][12];
       end
       11: begin
              muxOutConnector[0] = fifoOut[18][3];
              muxOutConnector[1] = fifoOut[19][3];
              muxOutConnector[2] = fifoOut[20][3];
              muxOutConnector[3] = fifoOut[21][3];
              muxOutConnector[4] = fifoOut[22][3];
              muxOutConnector[5] = fifoOut[23][3];
              muxOutConnector[6] = fifoOut[24][3];
              muxOutConnector[7] = fifoOut[26][10];
              muxOutConnector[8] = fifoOut[27][10];
              muxOutConnector[9] = fifoOut[28][10];
              muxOutConnector[10] = fifoOut[29][10];
              muxOutConnector[11] = fifoOut[30][10];
              muxOutConnector[12] = fifoOut[31][10];
              muxOutConnector[13] = fifoOut[32][10];
              muxOutConnector[14] = fifoOut[33][10];
              muxOutConnector[15] = fifoOut[34][10];
              muxOutConnector[16] = fifoOut[35][10];
              muxOutConnector[17] = fifoOut[36][10];
              muxOutConnector[18] = fifoOut[37][10];
              muxOutConnector[19] = fifoOut[38][10];
              muxOutConnector[20] = fifoOut[39][10];
              muxOutConnector[21] = fifoOut[40][10];
              muxOutConnector[22] = fifoOut[41][10];
              muxOutConnector[23] = fifoOut[42][10];
              muxOutConnector[24] = fifoOut[43][10];
              muxOutConnector[25] = fifoOut[44][10];
              muxOutConnector[26] = fifoOut[42][0];
              muxOutConnector[27] = fifoOut[43][0];
              muxOutConnector[28] = fifoOut[44][0];
              muxOutConnector[29] = fifoOut[45][0];
              muxOutConnector[30] = fifoOut[46][0];
              muxOutConnector[31] = fifoOut[47][0];
              muxOutConnector[32] = fifoOut[48][0];
              muxOutConnector[33] = fifoOut[49][0];
              muxOutConnector[34] = fifoOut[50][0];
              muxOutConnector[35] = fifoOut[51][0];
              muxOutConnector[36] = fifoOut[26][12];
              muxOutConnector[37] = fifoOut[27][12];
              muxOutConnector[38] = fifoOut[28][12];
              muxOutConnector[39] = fifoOut[29][12];
              muxOutConnector[40] = fifoOut[30][12];
              muxOutConnector[41] = fifoOut[31][12];
              muxOutConnector[42] = fifoOut[32][12];
              muxOutConnector[43] = fifoOut[33][12];
              muxOutConnector[44] = fifoOut[34][12];
              muxOutConnector[45] = fifoOut[35][12];
              muxOutConnector[46] = fifoOut[36][12];
              muxOutConnector[47] = fifoOut[37][12];
              muxOutConnector[48] = fifoOut[38][12];
              muxOutConnector[49] = fifoOut[39][12];
              muxOutConnector[50] = fifoOut[40][12];
              muxOutConnector[51] = fifoOut[41][12];
       end
       12: begin
              muxOutConnector[0] = fifoOut[45][11];
              muxOutConnector[1] = fifoOut[46][11];
              muxOutConnector[2] = fifoOut[47][11];
              muxOutConnector[3] = fifoOut[48][11];
              muxOutConnector[4] = fifoOut[49][11];
              muxOutConnector[5] = fifoOut[50][11];
              muxOutConnector[6] = fifoOut[51][11];
              muxOutConnector[7] = fifoOut[26][10];
              muxOutConnector[8] = fifoOut[27][10];
              muxOutConnector[9] = fifoOut[28][10];
              muxOutConnector[10] = fifoOut[29][10];
              muxOutConnector[11] = fifoOut[30][10];
              muxOutConnector[12] = fifoOut[31][10];
              muxOutConnector[13] = fifoOut[32][10];
              muxOutConnector[14] = fifoOut[33][10];
              muxOutConnector[15] = fifoOut[34][10];
              muxOutConnector[16] = fifoOut[35][10];
              muxOutConnector[17] = fifoOut[36][10];
              muxOutConnector[18] = fifoOut[37][10];
              muxOutConnector[19] = fifoOut[38][10];
              muxOutConnector[20] = fifoOut[39][10];
              muxOutConnector[21] = fifoOut[40][10];
              muxOutConnector[22] = fifoOut[41][10];
              muxOutConnector[23] = fifoOut[42][10];
              muxOutConnector[24] = fifoOut[43][10];
              muxOutConnector[25] = fifoOut[44][10];
              muxOutConnector[26] = fifoOut[42][0];
              muxOutConnector[27] = fifoOut[43][0];
              muxOutConnector[28] = fifoOut[0][11];
              muxOutConnector[29] = fifoOut[1][11];
              muxOutConnector[30] = fifoOut[2][11];
              muxOutConnector[31] = fifoOut[3][11];
              muxOutConnector[32] = fifoOut[4][11];
              muxOutConnector[33] = fifoOut[5][11];
              muxOutConnector[34] = fifoOut[6][11];
              muxOutConnector[35] = fifoOut[7][11];
              muxOutConnector[36] = fifoOut[26][12];
              muxOutConnector[37] = fifoOut[27][12];
              muxOutConnector[38] = fifoOut[28][12];
              muxOutConnector[39] = fifoOut[29][12];
              muxOutConnector[40] = fifoOut[30][12];
              muxOutConnector[41] = fifoOut[31][12];
              muxOutConnector[42] = fifoOut[32][12];
              muxOutConnector[43] = fifoOut[33][12];
              muxOutConnector[44] = fifoOut[34][12];
              muxOutConnector[45] = fifoOut[35][12];
              muxOutConnector[46] = fifoOut[36][12];
              muxOutConnector[47] = fifoOut[37][12];
              muxOutConnector[48] = fifoOut[38][12];
              muxOutConnector[49] = fifoOut[39][12];
              muxOutConnector[50] = fifoOut[40][12];
              muxOutConnector[51] = fifoOut[41][12];
       end
       13: begin
              muxOutConnector[0] = fifoOut[45][11];
              muxOutConnector[1] = fifoOut[46][11];
              muxOutConnector[2] = fifoOut[47][11];
              muxOutConnector[3] = fifoOut[48][11];
              muxOutConnector[4] = fifoOut[49][11];
              muxOutConnector[5] = fifoOut[50][11];
              muxOutConnector[6] = fifoOut[51][11];
              muxOutConnector[7] = fifoOut[26][10];
              muxOutConnector[8] = fifoOut[27][10];
              muxOutConnector[9] = fifoOut[28][10];
              muxOutConnector[10] = fifoOut[29][10];
              muxOutConnector[11] = fifoOut[30][10];
              muxOutConnector[12] = fifoOut[31][10];
              muxOutConnector[13] = fifoOut[32][10];
              muxOutConnector[14] = fifoOut[33][10];
              muxOutConnector[15] = fifoOut[34][10];
              muxOutConnector[16] = fifoOut[35][10];
              muxOutConnector[17] = fifoOut[36][10];
              muxOutConnector[18] = fifoOut[37][10];
              muxOutConnector[19] = fifoOut[38][10];
              muxOutConnector[20] = fifoOut[39][10];
              muxOutConnector[21] = fifoOut[40][10];
              muxOutConnector[22] = fifoOut[41][10];
              muxOutConnector[23] = fifoOut[42][10];
              muxOutConnector[24] = fifoOut[43][10];
              muxOutConnector[25] = fifoOut[44][10];
              muxOutConnector[26] = fifoOut[24][12];
              muxOutConnector[27] = fifoOut[25][12];
              muxOutConnector[28] = fifoOut[0][11];
              muxOutConnector[29] = fifoOut[1][11];
              muxOutConnector[30] = fifoOut[2][11];
              muxOutConnector[31] = fifoOut[3][11];
              muxOutConnector[32] = fifoOut[4][11];
              muxOutConnector[33] = fifoOut[5][11];
              muxOutConnector[34] = fifoOut[6][11];
              muxOutConnector[35] = fifoOut[7][11];
              muxOutConnector[36] = fifoOut[8][11];
              muxOutConnector[37] = fifoOut[9][11];
              muxOutConnector[38] = fifoOut[10][11];
              muxOutConnector[39] = fifoOut[11][11];
              muxOutConnector[40] = fifoOut[12][11];
              muxOutConnector[41] = fifoOut[13][11];
              muxOutConnector[42] = fifoOut[14][11];
              muxOutConnector[43] = fifoOut[15][11];
              muxOutConnector[44] = fifoOut[16][11];
              muxOutConnector[45] = fifoOut[17][11];
              muxOutConnector[46] = fifoOut[18][11];
              muxOutConnector[47] = fifoOut[19][11];
              muxOutConnector[48] = fifoOut[20][11];
              muxOutConnector[49] = fifoOut[21][11];
              muxOutConnector[50] = fifoOut[22][11];
              muxOutConnector[51] = fifoOut[23][11];
       end
       14: begin
              muxOutConnector[0] = fifoOut[45][11];
              muxOutConnector[1] = fifoOut[46][11];
              muxOutConnector[2] = fifoOut[47][11];
              muxOutConnector[3] = fifoOut[48][11];
              muxOutConnector[4] = fifoOut[49][11];
              muxOutConnector[5] = fifoOut[50][11];
              muxOutConnector[6] = fifoOut[51][11];
              muxOutConnector[7] = fifoOut[26][10];
              muxOutConnector[8] = fifoOut[27][10];
              muxOutConnector[9] = fifoOut[28][10];
              muxOutConnector[10] = fifoOut[29][10];
              muxOutConnector[11] = fifoOut[30][10];
              muxOutConnector[12] = fifoOut[31][10];
              muxOutConnector[13] = fifoOut[32][10];
              muxOutConnector[14] = fifoOut[33][10];
              muxOutConnector[15] = fifoOut[34][10];
              muxOutConnector[16] = fifoOut[35][10];
              muxOutConnector[17] = fifoOut[36][10];
              muxOutConnector[18] = fifoOut[37][10];
              muxOutConnector[19] = fifoOut[38][10];
              muxOutConnector[20] = fifoOut[39][10];
              muxOutConnector[21] = fifoOut[40][10];
              muxOutConnector[22] = fifoOut[41][10];
              muxOutConnector[23] = fifoOut[42][10];
              muxOutConnector[24] = fifoOut[43][10];
              muxOutConnector[25] = fifoOut[44][10];
              muxOutConnector[26] = fifoOut[24][12];
              muxOutConnector[27] = fifoOut[25][12];
              muxOutConnector[28] = fifoOut[0][11];
              muxOutConnector[29] = fifoOut[1][11];
              muxOutConnector[30] = fifoOut[2][11];
              muxOutConnector[31] = fifoOut[3][11];
              muxOutConnector[32] = fifoOut[4][11];
              muxOutConnector[33] = fifoOut[5][11];
              muxOutConnector[34] = fifoOut[6][11];
              muxOutConnector[35] = fifoOut[7][11];
              muxOutConnector[36] = fifoOut[8][11];
              muxOutConnector[37] = fifoOut[9][11];
              muxOutConnector[38] = fifoOut[10][11];
              muxOutConnector[39] = fifoOut[11][11];
              muxOutConnector[40] = fifoOut[12][11];
              muxOutConnector[41] = fifoOut[13][11];
              muxOutConnector[42] = fifoOut[14][11];
              muxOutConnector[43] = fifoOut[15][11];
              muxOutConnector[44] = fifoOut[16][11];
              muxOutConnector[45] = fifoOut[17][11];
              muxOutConnector[46] = fifoOut[18][11];
              muxOutConnector[47] = fifoOut[19][11];
              muxOutConnector[48] = fifoOut[20][11];
              muxOutConnector[49] = fifoOut[21][11];
              muxOutConnector[50] = fifoOut[22][11];
              muxOutConnector[51] = fifoOut[23][11];
       end
       15: begin
              muxOutConnector[0] = fifoOut[45][11];
              muxOutConnector[1] = fifoOut[46][11];
              muxOutConnector[2] = fifoOut[47][11];
              muxOutConnector[3] = fifoOut[48][11];
              muxOutConnector[4] = fifoOut[49][11];
              muxOutConnector[5] = fifoOut[50][11];
              muxOutConnector[6] = fifoOut[51][11];
              muxOutConnector[7] = fifoOut[26][10];
              muxOutConnector[8] = fifoOut[27][10];
              muxOutConnector[9] = fifoOut[28][10];
              muxOutConnector[10] = fifoOut[29][10];
              muxOutConnector[11] = fifoOut[30][10];
              muxOutConnector[12] = fifoOut[31][10];
              muxOutConnector[13] = fifoOut[32][10];
              muxOutConnector[14] = fifoOut[33][10];
              muxOutConnector[15] = fifoOut[34][10];
              muxOutConnector[16] = fifoOut[35][10];
              muxOutConnector[17] = fifoOut[36][10];
              muxOutConnector[18] = fifoOut[37][10];
              muxOutConnector[19] = fifoOut[38][10];
              muxOutConnector[20] = fifoOut[39][10];
              muxOutConnector[21] = fifoOut[40][10];
              muxOutConnector[22] = fifoOut[41][10];
              muxOutConnector[23] = fifoOut[42][10];
              muxOutConnector[24] = fifoOut[43][10];
              muxOutConnector[25] = fifoOut[44][10];
              muxOutConnector[26] = fifoOut[24][12];
              muxOutConnector[27] = fifoOut[25][12];
              muxOutConnector[28] = fifoOut[0][11];
              muxOutConnector[29] = fifoOut[1][11];
              muxOutConnector[30] = fifoOut[2][11];
              muxOutConnector[31] = fifoOut[3][11];
              muxOutConnector[32] = fifoOut[4][11];
              muxOutConnector[33] = fifoOut[5][11];
              muxOutConnector[34] = fifoOut[6][11];
              muxOutConnector[35] = fifoOut[7][11];
              muxOutConnector[36] = fifoOut[8][11];
              muxOutConnector[37] = fifoOut[9][11];
              muxOutConnector[38] = fifoOut[10][11];
              muxOutConnector[39] = fifoOut[11][11];
              muxOutConnector[40] = fifoOut[12][11];
              muxOutConnector[41] = fifoOut[13][11];
              muxOutConnector[42] = fifoOut[14][11];
              muxOutConnector[43] = fifoOut[15][11];
              muxOutConnector[44] = fifoOut[16][11];
              muxOutConnector[45] = fifoOut[17][11];
              muxOutConnector[46] = fifoOut[18][11];
              muxOutConnector[47] = fifoOut[19][11];
              muxOutConnector[48] = fifoOut[20][11];
              muxOutConnector[49] = fifoOut[21][11];
              muxOutConnector[50] = fifoOut[22][11];
              muxOutConnector[51] = fifoOut[23][11];
       end
       16: begin
              muxOutConnector[0] = fifoOut[45][11];
              muxOutConnector[1] = fifoOut[46][11];
              muxOutConnector[2] = fifoOut[47][11];
              muxOutConnector[3] = fifoOut[48][11];
              muxOutConnector[4] = fifoOut[49][11];
              muxOutConnector[5] = fifoOut[50][11];
              muxOutConnector[6] = fifoOut[51][11];
              muxOutConnector[7] = fifoOut[26][10];
              muxOutConnector[8] = fifoOut[27][10];
              muxOutConnector[9] = fifoOut[28][10];
              muxOutConnector[10] = fifoOut[29][10];
              muxOutConnector[11] = fifoOut[30][10];
              muxOutConnector[12] = fifoOut[31][10];
              muxOutConnector[13] = fifoOut[32][10];
              muxOutConnector[14] = fifoOut[33][10];
              muxOutConnector[15] = fifoOut[34][10];
              muxOutConnector[16] = fifoOut[35][10];
              muxOutConnector[17] = fifoOut[36][10];
              muxOutConnector[18] = fifoOut[37][10];
              muxOutConnector[19] = fifoOut[38][10];
              muxOutConnector[20] = fifoOut[39][10];
              muxOutConnector[21] = fifoOut[40][10];
              muxOutConnector[22] = fifoOut[41][10];
              muxOutConnector[23] = fifoOut[42][10];
              muxOutConnector[24] = fifoOut[43][10];
              muxOutConnector[25] = fifoOut[44][10];
              muxOutConnector[26] = fifoOut[24][12];
              muxOutConnector[27] = fifoOut[25][12];
              muxOutConnector[28] = fifoOut[0][11];
              muxOutConnector[29] = fifoOut[1][11];
              muxOutConnector[30] = fifoOut[2][11];
              muxOutConnector[31] = fifoOut[3][11];
              muxOutConnector[32] = fifoOut[4][11];
              muxOutConnector[33] = fifoOut[5][11];
              muxOutConnector[34] = fifoOut[6][11];
              muxOutConnector[35] = fifoOut[7][11];
              muxOutConnector[36] = fifoOut[8][11];
              muxOutConnector[37] = fifoOut[9][11];
              muxOutConnector[38] = fifoOut[10][11];
              muxOutConnector[39] = fifoOut[11][11];
              muxOutConnector[40] = fifoOut[12][11];
              muxOutConnector[41] = fifoOut[13][11];
              muxOutConnector[42] = fifoOut[14][11];
              muxOutConnector[43] = fifoOut[15][11];
              muxOutConnector[44] = fifoOut[16][11];
              muxOutConnector[45] = fifoOut[17][11];
              muxOutConnector[46] = fifoOut[18][11];
              muxOutConnector[47] = fifoOut[19][11];
              muxOutConnector[48] = fifoOut[20][11];
              muxOutConnector[49] = fifoOut[21][11];
              muxOutConnector[50] = fifoOut[22][11];
              muxOutConnector[51] = fifoOut[23][11];
       end
       17: begin
              muxOutConnector[0] = fifoOut[45][11];
              muxOutConnector[1] = fifoOut[46][11];
              muxOutConnector[2] = fifoOut[47][11];
              muxOutConnector[3] = fifoOut[48][11];
              muxOutConnector[4] = fifoOut[49][11];
              muxOutConnector[5] = fifoOut[50][11];
              muxOutConnector[6] = fifoOut[51][11];
              muxOutConnector[7] = fifoOut[26][10];
              muxOutConnector[8] = fifoOut[27][10];
              muxOutConnector[9] = fifoOut[28][10];
              muxOutConnector[10] = fifoOut[29][10];
              muxOutConnector[11] = fifoOut[30][10];
              muxOutConnector[12] = fifoOut[31][10];
              muxOutConnector[13] = fifoOut[32][10];
              muxOutConnector[14] = fifoOut[33][10];
              muxOutConnector[15] = fifoOut[34][10];
              muxOutConnector[16] = fifoOut[35][10];
              muxOutConnector[17] = fifoOut[36][10];
              muxOutConnector[18] = fifoOut[37][10];
              muxOutConnector[19] = fifoOut[38][10];
              muxOutConnector[20] = fifoOut[39][10];
              muxOutConnector[21] = fifoOut[40][10];
              muxOutConnector[22] = fifoOut[41][10];
              muxOutConnector[23] = fifoOut[42][10];
              muxOutConnector[24] = fifoOut[43][10];
              muxOutConnector[25] = fifoOut[44][10];
              muxOutConnector[26] = fifoOut[24][12];
              muxOutConnector[27] = fifoOut[25][12];
              muxOutConnector[28] = fifoOut[0][11];
              muxOutConnector[29] = fifoOut[1][11];
              muxOutConnector[30] = fifoOut[2][11];
              muxOutConnector[31] = fifoOut[3][11];
              muxOutConnector[32] = fifoOut[4][11];
              muxOutConnector[33] = fifoOut[5][11];
              muxOutConnector[34] = fifoOut[6][11];
              muxOutConnector[35] = fifoOut[7][11];
              muxOutConnector[36] = fifoOut[8][11];
              muxOutConnector[37] = fifoOut[9][11];
              muxOutConnector[38] = fifoOut[10][11];
              muxOutConnector[39] = fifoOut[11][11];
              muxOutConnector[40] = fifoOut[12][11];
              muxOutConnector[41] = fifoOut[13][11];
              muxOutConnector[42] = fifoOut[14][11];
              muxOutConnector[43] = fifoOut[15][11];
              muxOutConnector[44] = fifoOut[16][11];
              muxOutConnector[45] = fifoOut[17][11];
              muxOutConnector[46] = fifoOut[18][11];
              muxOutConnector[47] = fifoOut[19][11];
              muxOutConnector[48] = fifoOut[20][11];
              muxOutConnector[49] = fifoOut[21][11];
              muxOutConnector[50] = fifoOut[22][11];
              muxOutConnector[51] = fifoOut[23][11];
       end
       18: begin
              muxOutConnector[0] = fifoOut[45][11];
              muxOutConnector[1] = fifoOut[46][11];
              muxOutConnector[2] = fifoOut[47][11];
              muxOutConnector[3] = fifoOut[48][11];
              muxOutConnector[4] = fifoOut[49][11];
              muxOutConnector[5] = fifoOut[50][11];
              muxOutConnector[6] = fifoOut[51][11];
              muxOutConnector[7] = fifoOut[26][10];
              muxOutConnector[8] = fifoOut[27][10];
              muxOutConnector[9] = fifoOut[28][10];
              muxOutConnector[10] = fifoOut[29][10];
              muxOutConnector[11] = fifoOut[30][10];
              muxOutConnector[12] = fifoOut[31][10];
              muxOutConnector[13] = fifoOut[32][10];
              muxOutConnector[14] = fifoOut[33][10];
              muxOutConnector[15] = fifoOut[34][10];
              muxOutConnector[16] = fifoOut[35][10];
              muxOutConnector[17] = fifoOut[36][10];
              muxOutConnector[18] = fifoOut[37][10];
              muxOutConnector[19] = fifoOut[38][10];
              muxOutConnector[20] = fifoOut[39][10];
              muxOutConnector[21] = fifoOut[40][10];
              muxOutConnector[22] = fifoOut[41][10];
              muxOutConnector[23] = fifoOut[42][10];
              muxOutConnector[24] = fifoOut[43][10];
              muxOutConnector[25] = fifoOut[44][10];
              muxOutConnector[26] = fifoOut[24][12];
              muxOutConnector[27] = fifoOut[25][12];
              muxOutConnector[28] = fifoOut[0][11];
              muxOutConnector[29] = fifoOut[1][11];
              muxOutConnector[30] = fifoOut[2][11];
              muxOutConnector[31] = fifoOut[3][11];
              muxOutConnector[32] = fifoOut[4][11];
              muxOutConnector[33] = fifoOut[5][11];
              muxOutConnector[34] = fifoOut[6][11];
              muxOutConnector[35] = fifoOut[7][11];
              muxOutConnector[36] = fifoOut[8][11];
              muxOutConnector[37] = fifoOut[9][11];
              muxOutConnector[38] = fifoOut[10][11];
              muxOutConnector[39] = fifoOut[11][11];
              muxOutConnector[40] = fifoOut[12][11];
              muxOutConnector[41] = fifoOut[13][11];
              muxOutConnector[42] = fifoOut[14][11];
              muxOutConnector[43] = fifoOut[15][11];
              muxOutConnector[44] = fifoOut[16][11];
              muxOutConnector[45] = fifoOut[17][11];
              muxOutConnector[46] = fifoOut[18][11];
              muxOutConnector[47] = fifoOut[19][11];
              muxOutConnector[48] = fifoOut[20][11];
              muxOutConnector[49] = fifoOut[21][11];
              muxOutConnector[50] = fifoOut[22][11];
              muxOutConnector[51] = fifoOut[23][11];
       end
       19: begin
              muxOutConnector[0] = fifoOut[45][11];
              muxOutConnector[1] = fifoOut[46][11];
              muxOutConnector[2] = fifoOut[47][11];
              muxOutConnector[3] = fifoOut[48][11];
              muxOutConnector[4] = fifoOut[49][11];
              muxOutConnector[5] = fifoOut[50][11];
              muxOutConnector[6] = fifoOut[51][11];
              muxOutConnector[7] = fifoOut[26][10];
              muxOutConnector[8] = fifoOut[27][10];
              muxOutConnector[9] = fifoOut[28][10];
              muxOutConnector[10] = fifoOut[29][10];
              muxOutConnector[11] = fifoOut[30][10];
              muxOutConnector[12] = fifoOut[31][10];
              muxOutConnector[13] = fifoOut[32][10];
              muxOutConnector[14] = fifoOut[33][10];
              muxOutConnector[15] = fifoOut[34][10];
              muxOutConnector[16] = fifoOut[35][10];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[24][12];
              muxOutConnector[27] = fifoOut[25][12];
              muxOutConnector[28] = fifoOut[0][11];
              muxOutConnector[29] = fifoOut[1][11];
              muxOutConnector[30] = fifoOut[2][11];
              muxOutConnector[31] = fifoOut[3][11];
              muxOutConnector[32] = fifoOut[4][11];
              muxOutConnector[33] = fifoOut[5][11];
              muxOutConnector[34] = fifoOut[6][11];
              muxOutConnector[35] = fifoOut[7][11];
              muxOutConnector[36] = fifoOut[8][11];
              muxOutConnector[37] = fifoOut[9][11];
              muxOutConnector[38] = fifoOut[10][11];
              muxOutConnector[39] = fifoOut[11][11];
              muxOutConnector[40] = fifoOut[12][11];
              muxOutConnector[41] = fifoOut[13][11];
              muxOutConnector[42] = fifoOut[14][11];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
