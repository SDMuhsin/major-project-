`timescale 1ns / 1ps
module LMem1To0_511_circ2_ys_yu_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 11;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input [ADDRESSWIDTH-1:0]unloadAddress;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            fifoOut[i][0] <= ly0InConnector[i];
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
       0: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = fifoOut[1][7][w-1];
              unloadMuxOut[31] = fifoOut[2][7][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[3][7][w-1];
              unloadMuxOut[1] = fifoOut[4][7][w-1];
              unloadMuxOut[2] = fifoOut[5][7][w-1];
              unloadMuxOut[3] = fifoOut[6][7][w-1];
              unloadMuxOut[4] = fifoOut[7][7][w-1];
              unloadMuxOut[5] = fifoOut[8][7][w-1];
              unloadMuxOut[6] = fifoOut[9][7][w-1];
              unloadMuxOut[7] = fifoOut[10][7][w-1];
              unloadMuxOut[8] = fifoOut[11][7][w-1];
              unloadMuxOut[9] = fifoOut[12][7][w-1];
              unloadMuxOut[10] = fifoOut[13][7][w-1];
              unloadMuxOut[11] = fifoOut[14][7][w-1];
              unloadMuxOut[12] = fifoOut[15][7][w-1];
              unloadMuxOut[13] = fifoOut[16][7][w-1];
              unloadMuxOut[14] = fifoOut[17][7][w-1];
              unloadMuxOut[15] = fifoOut[18][7][w-1];
              unloadMuxOut[16] = fifoOut[19][7][w-1];
              unloadMuxOut[17] = fifoOut[20][7][w-1];
              unloadMuxOut[18] = fifoOut[21][7][w-1];
              unloadMuxOut[19] = fifoOut[22][7][w-1];
              unloadMuxOut[20] = fifoOut[23][7][w-1];
              unloadMuxOut[21] = fifoOut[24][7][w-1];
              unloadMuxOut[22] = fifoOut[25][7][w-1];
              unloadMuxOut[23] = fifoOut[0][6][w-1];
              unloadMuxOut[24] = fifoOut[1][6][w-1];
              unloadMuxOut[25] = fifoOut[2][6][w-1];
              unloadMuxOut[26] = fifoOut[3][6][w-1];
              unloadMuxOut[27] = fifoOut[4][6][w-1];
              unloadMuxOut[28] = fifoOut[5][6][w-1];
              unloadMuxOut[29] = fifoOut[6][6][w-1];
              unloadMuxOut[30] = fifoOut[7][6][w-1];
              unloadMuxOut[31] = fifoOut[8][6][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[9][6][w-1];
              unloadMuxOut[1] = fifoOut[10][6][w-1];
              unloadMuxOut[2] = fifoOut[11][6][w-1];
              unloadMuxOut[3] = fifoOut[12][6][w-1];
              unloadMuxOut[4] = fifoOut[13][6][w-1];
              unloadMuxOut[5] = fifoOut[14][6][w-1];
              unloadMuxOut[6] = fifoOut[15][6][w-1];
              unloadMuxOut[7] = fifoOut[16][6][w-1];
              unloadMuxOut[8] = fifoOut[17][6][w-1];
              unloadMuxOut[9] = fifoOut[18][6][w-1];
              unloadMuxOut[10] = fifoOut[19][6][w-1];
              unloadMuxOut[11] = fifoOut[20][6][w-1];
              unloadMuxOut[12] = fifoOut[21][6][w-1];
              unloadMuxOut[13] = fifoOut[22][6][w-1];
              unloadMuxOut[14] = fifoOut[23][6][w-1];
              unloadMuxOut[15] = fifoOut[24][6][w-1];
              unloadMuxOut[16] = fifoOut[25][6][w-1];
              unloadMuxOut[17] = fifoOut[0][5][w-1];
              unloadMuxOut[18] = fifoOut[1][5][w-1];
              unloadMuxOut[19] = fifoOut[2][5][w-1];
              unloadMuxOut[20] = fifoOut[3][5][w-1];
              unloadMuxOut[21] = fifoOut[4][5][w-1];
              unloadMuxOut[22] = fifoOut[5][5][w-1];
              unloadMuxOut[23] = fifoOut[6][5][w-1];
              unloadMuxOut[24] = fifoOut[7][5][w-1];
              unloadMuxOut[25] = fifoOut[8][5][w-1];
              unloadMuxOut[26] = fifoOut[9][5][w-1];
              unloadMuxOut[27] = fifoOut[10][5][w-1];
              unloadMuxOut[28] = fifoOut[11][5][w-1];
              unloadMuxOut[29] = fifoOut[12][5][w-1];
              unloadMuxOut[30] = fifoOut[13][5][w-1];
              unloadMuxOut[31] = fifoOut[14][5][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[15][5][w-1];
              unloadMuxOut[1] = fifoOut[16][5][w-1];
              unloadMuxOut[2] = fifoOut[17][5][w-1];
              unloadMuxOut[3] = fifoOut[18][5][w-1];
              unloadMuxOut[4] = fifoOut[19][5][w-1];
              unloadMuxOut[5] = fifoOut[20][5][w-1];
              unloadMuxOut[6] = fifoOut[21][5][w-1];
              unloadMuxOut[7] = fifoOut[22][5][w-1];
              unloadMuxOut[8] = fifoOut[23][5][w-1];
              unloadMuxOut[9] = fifoOut[24][5][w-1];
              unloadMuxOut[10] = fifoOut[25][5][w-1];
              unloadMuxOut[11] = fifoOut[0][4][w-1];
              unloadMuxOut[12] = fifoOut[1][4][w-1];
              unloadMuxOut[13] = fifoOut[2][4][w-1];
              unloadMuxOut[14] = fifoOut[3][4][w-1];
              unloadMuxOut[15] = fifoOut[4][4][w-1];
              unloadMuxOut[16] = fifoOut[5][4][w-1];
              unloadMuxOut[17] = fifoOut[6][4][w-1];
              unloadMuxOut[18] = fifoOut[7][4][w-1];
              unloadMuxOut[19] = fifoOut[8][4][w-1];
              unloadMuxOut[20] = fifoOut[9][4][w-1];
              unloadMuxOut[21] = fifoOut[10][4][w-1];
              unloadMuxOut[22] = fifoOut[11][4][w-1];
              unloadMuxOut[23] = fifoOut[12][4][w-1];
              unloadMuxOut[24] = fifoOut[13][4][w-1];
              unloadMuxOut[25] = fifoOut[14][4][w-1];
              unloadMuxOut[26] = fifoOut[15][4][w-1];
              unloadMuxOut[27] = fifoOut[16][4][w-1];
              unloadMuxOut[28] = fifoOut[17][4][w-1];
              unloadMuxOut[29] = fifoOut[18][4][w-1];
              unloadMuxOut[30] = fifoOut[19][4][w-1];
              unloadMuxOut[31] = fifoOut[20][4][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[21][4][w-1];
              unloadMuxOut[1] = fifoOut[22][4][w-1];
              unloadMuxOut[2] = fifoOut[23][4][w-1];
              unloadMuxOut[3] = fifoOut[24][4][w-1];
              unloadMuxOut[4] = fifoOut[25][4][w-1];
              unloadMuxOut[5] = fifoOut[0][3][w-1];
              unloadMuxOut[6] = fifoOut[1][3][w-1];
              unloadMuxOut[7] = fifoOut[2][3][w-1];
              unloadMuxOut[8] = fifoOut[3][3][w-1];
              unloadMuxOut[9] = fifoOut[4][3][w-1];
              unloadMuxOut[10] = fifoOut[5][3][w-1];
              unloadMuxOut[11] = fifoOut[6][3][w-1];
              unloadMuxOut[12] = fifoOut[7][3][w-1];
              unloadMuxOut[13] = fifoOut[8][3][w-1];
              unloadMuxOut[14] = fifoOut[9][3][w-1];
              unloadMuxOut[15] = fifoOut[10][3][w-1];
              unloadMuxOut[16] = fifoOut[11][3][w-1];
              unloadMuxOut[17] = fifoOut[12][3][w-1];
              unloadMuxOut[18] = fifoOut[13][3][w-1];
              unloadMuxOut[19] = fifoOut[14][3][w-1];
              unloadMuxOut[20] = fifoOut[15][3][w-1];
              unloadMuxOut[21] = fifoOut[16][3][w-1];
              unloadMuxOut[22] = fifoOut[17][3][w-1];
              unloadMuxOut[23] = fifoOut[18][3][w-1];
              unloadMuxOut[24] = fifoOut[19][3][w-1];
              unloadMuxOut[25] = fifoOut[20][3][w-1];
              unloadMuxOut[26] = fifoOut[21][3][w-1];
              unloadMuxOut[27] = fifoOut[22][3][w-1];
              unloadMuxOut[28] = fifoOut[23][3][w-1];
              unloadMuxOut[29] = fifoOut[24][3][w-1];
              unloadMuxOut[30] = fifoOut[25][3][w-1];
              unloadMuxOut[31] = fifoOut[0][2][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[1][2][w-1];
              unloadMuxOut[1] = fifoOut[2][2][w-1];
              unloadMuxOut[2] = fifoOut[3][2][w-1];
              unloadMuxOut[3] = fifoOut[4][2][w-1];
              unloadMuxOut[4] = fifoOut[5][2][w-1];
              unloadMuxOut[5] = fifoOut[6][2][w-1];
              unloadMuxOut[6] = fifoOut[7][2][w-1];
              unloadMuxOut[7] = fifoOut[8][2][w-1];
              unloadMuxOut[8] = fifoOut[9][2][w-1];
              unloadMuxOut[9] = fifoOut[10][2][w-1];
              unloadMuxOut[10] = fifoOut[11][2][w-1];
              unloadMuxOut[11] = fifoOut[12][2][w-1];
              unloadMuxOut[12] = fifoOut[13][2][w-1];
              unloadMuxOut[13] = fifoOut[14][2][w-1];
              unloadMuxOut[14] = fifoOut[15][2][w-1];
              unloadMuxOut[15] = fifoOut[16][2][w-1];
              unloadMuxOut[16] = fifoOut[17][2][w-1];
              unloadMuxOut[17] = fifoOut[18][2][w-1];
              unloadMuxOut[18] = fifoOut[19][2][w-1];
              unloadMuxOut[19] = fifoOut[20][2][w-1];
              unloadMuxOut[20] = fifoOut[21][2][w-1];
              unloadMuxOut[21] = fifoOut[22][2][w-1];
              unloadMuxOut[22] = fifoOut[23][2][w-1];
              unloadMuxOut[23] = fifoOut[24][2][w-1];
              unloadMuxOut[24] = fifoOut[25][2][w-1];
              unloadMuxOut[25] = fifoOut[0][1][w-1];
              unloadMuxOut[26] = fifoOut[1][1][w-1];
              unloadMuxOut[27] = fifoOut[2][1][w-1];
              unloadMuxOut[28] = fifoOut[26][10][w-1];
              unloadMuxOut[29] = fifoOut[27][10][w-1];
              unloadMuxOut[30] = fifoOut[28][10][w-1];
              unloadMuxOut[31] = fifoOut[29][10][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[30][10][w-1];
              unloadMuxOut[1] = fifoOut[31][10][w-1];
              unloadMuxOut[2] = fifoOut[32][10][w-1];
              unloadMuxOut[3] = fifoOut[33][10][w-1];
              unloadMuxOut[4] = fifoOut[34][10][w-1];
              unloadMuxOut[5] = fifoOut[35][10][w-1];
              unloadMuxOut[6] = fifoOut[36][10][w-1];
              unloadMuxOut[7] = fifoOut[37][10][w-1];
              unloadMuxOut[8] = fifoOut[38][10][w-1];
              unloadMuxOut[9] = fifoOut[39][10][w-1];
              unloadMuxOut[10] = fifoOut[40][10][w-1];
              unloadMuxOut[11] = fifoOut[41][10][w-1];
              unloadMuxOut[12] = fifoOut[42][10][w-1];
              unloadMuxOut[13] = fifoOut[43][10][w-1];
              unloadMuxOut[14] = fifoOut[44][10][w-1];
              unloadMuxOut[15] = fifoOut[45][10][w-1];
              unloadMuxOut[16] = fifoOut[46][10][w-1];
              unloadMuxOut[17] = fifoOut[47][10][w-1];
              unloadMuxOut[18] = fifoOut[48][10][w-1];
              unloadMuxOut[19] = fifoOut[49][10][w-1];
              unloadMuxOut[20] = fifoOut[50][10][w-1];
              unloadMuxOut[21] = fifoOut[51][10][w-1];
              unloadMuxOut[22] = fifoOut[26][9][w-1];
              unloadMuxOut[23] = fifoOut[27][9][w-1];
              unloadMuxOut[24] = fifoOut[28][9][w-1];
              unloadMuxOut[25] = fifoOut[29][9][w-1];
              unloadMuxOut[26] = fifoOut[30][9][w-1];
              unloadMuxOut[27] = fifoOut[31][9][w-1];
              unloadMuxOut[28] = fifoOut[32][9][w-1];
              unloadMuxOut[29] = fifoOut[33][9][w-1];
              unloadMuxOut[30] = fifoOut[34][9][w-1];
              unloadMuxOut[31] = fifoOut[35][9][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[36][9][w-1];
              unloadMuxOut[1] = fifoOut[37][9][w-1];
              unloadMuxOut[2] = fifoOut[38][9][w-1];
              unloadMuxOut[3] = fifoOut[39][9][w-1];
              unloadMuxOut[4] = fifoOut[40][9][w-1];
              unloadMuxOut[5] = fifoOut[41][9][w-1];
              unloadMuxOut[6] = fifoOut[42][9][w-1];
              unloadMuxOut[7] = fifoOut[43][9][w-1];
              unloadMuxOut[8] = fifoOut[44][9][w-1];
              unloadMuxOut[9] = fifoOut[45][9][w-1];
              unloadMuxOut[10] = fifoOut[46][9][w-1];
              unloadMuxOut[11] = fifoOut[47][9][w-1];
              unloadMuxOut[12] = fifoOut[48][9][w-1];
              unloadMuxOut[13] = fifoOut[49][9][w-1];
              unloadMuxOut[14] = fifoOut[50][9][w-1];
              unloadMuxOut[15] = fifoOut[51][9][w-1];
              unloadMuxOut[16] = fifoOut[26][8][w-1];
              unloadMuxOut[17] = fifoOut[27][8][w-1];
              unloadMuxOut[18] = fifoOut[28][8][w-1];
              unloadMuxOut[19] = fifoOut[29][8][w-1];
              unloadMuxOut[20] = fifoOut[30][8][w-1];
              unloadMuxOut[21] = fifoOut[31][8][w-1];
              unloadMuxOut[22] = fifoOut[32][8][w-1];
              unloadMuxOut[23] = fifoOut[33][8][w-1];
              unloadMuxOut[24] = fifoOut[34][8][w-1];
              unloadMuxOut[25] = fifoOut[35][8][w-1];
              unloadMuxOut[26] = fifoOut[36][8][w-1];
              unloadMuxOut[27] = fifoOut[37][8][w-1];
              unloadMuxOut[28] = fifoOut[38][8][w-1];
              unloadMuxOut[29] = fifoOut[39][8][w-1];
              unloadMuxOut[30] = fifoOut[40][8][w-1];
              unloadMuxOut[31] = fifoOut[41][8][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[42][8][w-1];
              unloadMuxOut[1] = fifoOut[43][8][w-1];
              unloadMuxOut[2] = fifoOut[44][8][w-1];
              unloadMuxOut[3] = fifoOut[45][8][w-1];
              unloadMuxOut[4] = fifoOut[46][8][w-1];
              unloadMuxOut[5] = fifoOut[47][8][w-1];
              unloadMuxOut[6] = fifoOut[48][8][w-1];
              unloadMuxOut[7] = fifoOut[49][8][w-1];
              unloadMuxOut[8] = fifoOut[50][8][w-1];
              unloadMuxOut[9] = fifoOut[51][8][w-1];
              unloadMuxOut[10] = fifoOut[26][7][w-1];
              unloadMuxOut[11] = fifoOut[27][7][w-1];
              unloadMuxOut[12] = fifoOut[28][7][w-1];
              unloadMuxOut[13] = fifoOut[29][7][w-1];
              unloadMuxOut[14] = fifoOut[30][7][w-1];
              unloadMuxOut[15] = fifoOut[31][7][w-1];
              unloadMuxOut[16] = fifoOut[32][7][w-1];
              unloadMuxOut[17] = fifoOut[33][7][w-1];
              unloadMuxOut[18] = fifoOut[34][7][w-1];
              unloadMuxOut[19] = fifoOut[35][7][w-1];
              unloadMuxOut[20] = fifoOut[36][7][w-1];
              unloadMuxOut[21] = fifoOut[37][7][w-1];
              unloadMuxOut[22] = fifoOut[38][7][w-1];
              unloadMuxOut[23] = fifoOut[39][7][w-1];
              unloadMuxOut[24] = fifoOut[40][7][w-1];
              unloadMuxOut[25] = fifoOut[41][7][w-1];
              unloadMuxOut[26] = fifoOut[42][7][w-1];
              unloadMuxOut[27] = fifoOut[43][7][w-1];
              unloadMuxOut[28] = fifoOut[44][7][w-1];
              unloadMuxOut[29] = fifoOut[45][7][w-1];
              unloadMuxOut[30] = fifoOut[46][7][w-1];
              unloadMuxOut[31] = fifoOut[47][7][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[48][7][w-1];
              unloadMuxOut[1] = fifoOut[49][7][w-1];
              unloadMuxOut[2] = fifoOut[50][7][w-1];
              unloadMuxOut[3] = fifoOut[51][7][w-1];
              unloadMuxOut[4] = fifoOut[26][6][w-1];
              unloadMuxOut[5] = fifoOut[27][6][w-1];
              unloadMuxOut[6] = fifoOut[28][6][w-1];
              unloadMuxOut[7] = fifoOut[29][6][w-1];
              unloadMuxOut[8] = fifoOut[30][6][w-1];
              unloadMuxOut[9] = fifoOut[31][6][w-1];
              unloadMuxOut[10] = fifoOut[32][6][w-1];
              unloadMuxOut[11] = fifoOut[33][6][w-1];
              unloadMuxOut[12] = fifoOut[34][6][w-1];
              unloadMuxOut[13] = fifoOut[35][6][w-1];
              unloadMuxOut[14] = fifoOut[36][6][w-1];
              unloadMuxOut[15] = fifoOut[37][6][w-1];
              unloadMuxOut[16] = fifoOut[38][6][w-1];
              unloadMuxOut[17] = fifoOut[39][6][w-1];
              unloadMuxOut[18] = fifoOut[40][6][w-1];
              unloadMuxOut[19] = fifoOut[41][6][w-1];
              unloadMuxOut[20] = fifoOut[42][6][w-1];
              unloadMuxOut[21] = fifoOut[43][6][w-1];
              unloadMuxOut[22] = fifoOut[44][6][w-1];
              unloadMuxOut[23] = fifoOut[45][6][w-1];
              unloadMuxOut[24] = fifoOut[46][6][w-1];
              unloadMuxOut[25] = fifoOut[47][6][w-1];
              unloadMuxOut[26] = fifoOut[48][6][w-1];
              unloadMuxOut[27] = fifoOut[49][6][w-1];
              unloadMuxOut[28] = fifoOut[50][6][w-1];
              unloadMuxOut[29] = fifoOut[51][6][w-1];
              unloadMuxOut[30] = fifoOut[26][5][w-1];
              unloadMuxOut[31] = fifoOut[27][5][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[28][5][w-1];
              unloadMuxOut[1] = fifoOut[29][5][w-1];
              unloadMuxOut[2] = fifoOut[30][5][w-1];
              unloadMuxOut[3] = fifoOut[31][5][w-1];
              unloadMuxOut[4] = fifoOut[32][5][w-1];
              unloadMuxOut[5] = fifoOut[33][5][w-1];
              unloadMuxOut[6] = fifoOut[34][5][w-1];
              unloadMuxOut[7] = fifoOut[35][5][w-1];
              unloadMuxOut[8] = fifoOut[36][5][w-1];
              unloadMuxOut[9] = fifoOut[37][5][w-1];
              unloadMuxOut[10] = fifoOut[38][5][w-1];
              unloadMuxOut[11] = fifoOut[39][5][w-1];
              unloadMuxOut[12] = fifoOut[40][5][w-1];
              unloadMuxOut[13] = fifoOut[41][5][w-1];
              unloadMuxOut[14] = fifoOut[42][5][w-1];
              unloadMuxOut[15] = fifoOut[43][5][w-1];
              unloadMuxOut[16] = fifoOut[44][5][w-1];
              unloadMuxOut[17] = fifoOut[45][5][w-1];
              unloadMuxOut[18] = fifoOut[46][5][w-1];
              unloadMuxOut[19] = fifoOut[47][5][w-1];
              unloadMuxOut[20] = fifoOut[48][5][w-1];
              unloadMuxOut[21] = fifoOut[49][5][w-1];
              unloadMuxOut[22] = fifoOut[50][5][w-1];
              unloadMuxOut[23] = fifoOut[51][5][w-1];
              unloadMuxOut[24] = fifoOut[26][4][w-1];
              unloadMuxOut[25] = fifoOut[27][4][w-1];
              unloadMuxOut[26] = fifoOut[28][4][w-1];
              unloadMuxOut[27] = fifoOut[29][4][w-1];
              unloadMuxOut[28] = fifoOut[30][4][w-1];
              unloadMuxOut[29] = fifoOut[31][4][w-1];
              unloadMuxOut[30] = fifoOut[32][4][w-1];
              unloadMuxOut[31] = fifoOut[33][4][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[34][4][w-1];
              unloadMuxOut[1] = fifoOut[35][4][w-1];
              unloadMuxOut[2] = fifoOut[36][4][w-1];
              unloadMuxOut[3] = fifoOut[37][4][w-1];
              unloadMuxOut[4] = fifoOut[38][4][w-1];
              unloadMuxOut[5] = fifoOut[39][4][w-1];
              unloadMuxOut[6] = fifoOut[40][4][w-1];
              unloadMuxOut[7] = fifoOut[41][4][w-1];
              unloadMuxOut[8] = fifoOut[42][4][w-1];
              unloadMuxOut[9] = fifoOut[43][4][w-1];
              unloadMuxOut[10] = fifoOut[44][4][w-1];
              unloadMuxOut[11] = fifoOut[45][4][w-1];
              unloadMuxOut[12] = fifoOut[46][4][w-1];
              unloadMuxOut[13] = fifoOut[47][4][w-1];
              unloadMuxOut[14] = fifoOut[48][4][w-1];
              unloadMuxOut[15] = fifoOut[49][4][w-1];
              unloadMuxOut[16] = fifoOut[50][4][w-1];
              unloadMuxOut[17] = fifoOut[51][4][w-1];
              unloadMuxOut[18] = fifoOut[26][3][w-1];
              unloadMuxOut[19] = fifoOut[27][3][w-1];
              unloadMuxOut[20] = fifoOut[28][3][w-1];
              unloadMuxOut[21] = fifoOut[29][3][w-1];
              unloadMuxOut[22] = fifoOut[30][3][w-1];
              unloadMuxOut[23] = fifoOut[31][3][w-1];
              unloadMuxOut[24] = fifoOut[32][3][w-1];
              unloadMuxOut[25] = fifoOut[33][3][w-1];
              unloadMuxOut[26] = fifoOut[34][3][w-1];
              unloadMuxOut[27] = fifoOut[35][3][w-1];
              unloadMuxOut[28] = fifoOut[36][3][w-1];
              unloadMuxOut[29] = fifoOut[37][3][w-1];
              unloadMuxOut[30] = fifoOut[38][3][w-1];
              unloadMuxOut[31] = fifoOut[39][3][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[40][3][w-1];
              unloadMuxOut[1] = fifoOut[41][3][w-1];
              unloadMuxOut[2] = fifoOut[42][3][w-1];
              unloadMuxOut[3] = fifoOut[43][3][w-1];
              unloadMuxOut[4] = fifoOut[44][3][w-1];
              unloadMuxOut[5] = fifoOut[45][3][w-1];
              unloadMuxOut[6] = fifoOut[46][3][w-1];
              unloadMuxOut[7] = fifoOut[47][3][w-1];
              unloadMuxOut[8] = fifoOut[48][3][w-1];
              unloadMuxOut[9] = fifoOut[49][3][w-1];
              unloadMuxOut[10] = fifoOut[50][3][w-1];
              unloadMuxOut[11] = fifoOut[51][3][w-1];
              unloadMuxOut[12] = fifoOut[26][2][w-1];
              unloadMuxOut[13] = fifoOut[27][2][w-1];
              unloadMuxOut[14] = fifoOut[28][2][w-1];
              unloadMuxOut[15] = fifoOut[29][2][w-1];
              unloadMuxOut[16] = fifoOut[30][2][w-1];
              unloadMuxOut[17] = fifoOut[31][2][w-1];
              unloadMuxOut[18] = fifoOut[32][2][w-1];
              unloadMuxOut[19] = fifoOut[33][2][w-1];
              unloadMuxOut[20] = fifoOut[34][2][w-1];
              unloadMuxOut[21] = fifoOut[35][2][w-1];
              unloadMuxOut[22] = fifoOut[36][2][w-1];
              unloadMuxOut[23] = fifoOut[37][2][w-1];
              unloadMuxOut[24] = fifoOut[38][2][w-1];
              unloadMuxOut[25] = fifoOut[39][2][w-1];
              unloadMuxOut[26] = fifoOut[40][2][w-1];
              unloadMuxOut[27] = fifoOut[41][2][w-1];
              unloadMuxOut[28] = fifoOut[42][2][w-1];
              unloadMuxOut[29] = fifoOut[43][2][w-1];
              unloadMuxOut[30] = fifoOut[44][2][w-1];
              unloadMuxOut[31] = fifoOut[45][2][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[46][2][w-1];
              unloadMuxOut[1] = fifoOut[47][2][w-1];
              unloadMuxOut[2] = fifoOut[48][2][w-1];
              unloadMuxOut[3] = fifoOut[49][2][w-1];
              unloadMuxOut[4] = fifoOut[50][2][w-1];
              unloadMuxOut[5] = fifoOut[51][2][w-1];
              unloadMuxOut[6] = fifoOut[26][1][w-1];
              unloadMuxOut[7] = fifoOut[27][1][w-1];
              unloadMuxOut[8] = fifoOut[28][1][w-1];
              unloadMuxOut[9] = fifoOut[29][1][w-1];
              unloadMuxOut[10] = fifoOut[30][1][w-1];
              unloadMuxOut[11] = fifoOut[31][1][w-1];
              unloadMuxOut[12] = fifoOut[32][1][w-1];
              unloadMuxOut[13] = fifoOut[33][1][w-1];
              unloadMuxOut[14] = fifoOut[34][1][w-1];
              unloadMuxOut[15] = fifoOut[35][1][w-1];
              unloadMuxOut[16] = fifoOut[36][1][w-1];
              unloadMuxOut[17] = fifoOut[37][1][w-1];
              unloadMuxOut[18] = fifoOut[38][1][w-1];
              unloadMuxOut[19] = fifoOut[39][1][w-1];
              unloadMuxOut[20] = fifoOut[40][1][w-1];
              unloadMuxOut[21] = fifoOut[41][1][w-1];
              unloadMuxOut[22] = fifoOut[42][1][w-1];
              unloadMuxOut[23] = fifoOut[43][1][w-1];
              unloadMuxOut[24] = fifoOut[44][1][w-1];
              unloadMuxOut[25] = fifoOut[45][1][w-1];
              unloadMuxOut[26] = fifoOut[46][1][w-1];
              unloadMuxOut[27] = fifoOut[47][1][w-1];
              unloadMuxOut[28] = fifoOut[48][1][w-1];
              unloadMuxOut[29] = fifoOut[49][1][w-1];
              unloadMuxOut[30] = fifoOut[50][1][w-1];
              unloadMuxOut[31] = fifoOut[51][1][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[26][0][w-1];
              unloadMuxOut[1] = fifoOut[27][0][w-1];
              unloadMuxOut[2] = fifoOut[28][0][w-1];
              unloadMuxOut[3] = fifoOut[29][0][w-1];
              unloadMuxOut[4] = fifoOut[30][0][w-1];
              unloadMuxOut[5] = fifoOut[31][0][w-1];
              unloadMuxOut[6] = fifoOut[32][0][w-1];
              unloadMuxOut[7] = fifoOut[33][0][w-1];
              unloadMuxOut[8] = fifoOut[34][0][w-1];
              unloadMuxOut[9] = fifoOut[35][0][w-1];
              unloadMuxOut[10] = fifoOut[36][0][w-1];
              unloadMuxOut[11] = fifoOut[37][0][w-1];
              unloadMuxOut[12] = fifoOut[38][0][w-1];
              unloadMuxOut[13] = fifoOut[39][0][w-1];
              unloadMuxOut[14] = fifoOut[0][10][w-1];
              unloadMuxOut[15] = fifoOut[1][10][w-1];
              unloadMuxOut[16] = fifoOut[2][10][w-1];
              unloadMuxOut[17] = fifoOut[3][10][w-1];
              unloadMuxOut[18] = fifoOut[4][10][w-1];
              unloadMuxOut[19] = fifoOut[5][10][w-1];
              unloadMuxOut[20] = fifoOut[6][10][w-1];
              unloadMuxOut[21] = fifoOut[7][10][w-1];
              unloadMuxOut[22] = fifoOut[8][10][w-1];
              unloadMuxOut[23] = fifoOut[9][10][w-1];
              unloadMuxOut[24] = fifoOut[10][10][w-1];
              unloadMuxOut[25] = fifoOut[11][10][w-1];
              unloadMuxOut[26] = fifoOut[12][10][w-1];
              unloadMuxOut[27] = fifoOut[13][10][w-1];
              unloadMuxOut[28] = fifoOut[14][10][w-1];
              unloadMuxOut[29] = fifoOut[15][10][w-1];
              unloadMuxOut[30] = fifoOut[16][10][w-1];
              unloadMuxOut[31] = fifoOut[17][10][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[18][10][w-1];
              unloadMuxOut[1] = fifoOut[19][10][w-1];
              unloadMuxOut[2] = fifoOut[20][10][w-1];
              unloadMuxOut[3] = fifoOut[21][10][w-1];
              unloadMuxOut[4] = fifoOut[22][10][w-1];
              unloadMuxOut[5] = fifoOut[23][10][w-1];
              unloadMuxOut[6] = fifoOut[24][10][w-1];
              unloadMuxOut[7] = fifoOut[25][10][w-1];
              unloadMuxOut[8] = fifoOut[0][9][w-1];
              unloadMuxOut[9] = fifoOut[1][9][w-1];
              unloadMuxOut[10] = fifoOut[2][9][w-1];
              unloadMuxOut[11] = fifoOut[3][9][w-1];
              unloadMuxOut[12] = fifoOut[4][9][w-1];
              unloadMuxOut[13] = fifoOut[5][9][w-1];
              unloadMuxOut[14] = fifoOut[6][9][w-1];
              unloadMuxOut[15] = fifoOut[7][9][w-1];
              unloadMuxOut[16] = fifoOut[8][9][w-1];
              unloadMuxOut[17] = fifoOut[9][9][w-1];
              unloadMuxOut[18] = fifoOut[10][9][w-1];
              unloadMuxOut[19] = fifoOut[11][9][w-1];
              unloadMuxOut[20] = fifoOut[12][9][w-1];
              unloadMuxOut[21] = fifoOut[13][9][w-1];
              unloadMuxOut[22] = fifoOut[14][9][w-1];
              unloadMuxOut[23] = fifoOut[15][9][w-1];
              unloadMuxOut[24] = fifoOut[16][9][w-1];
              unloadMuxOut[25] = fifoOut[17][9][w-1];
              unloadMuxOut[26] = fifoOut[18][9][w-1];
              unloadMuxOut[27] = fifoOut[19][9][w-1];
              unloadMuxOut[28] = fifoOut[20][9][w-1];
              unloadMuxOut[29] = fifoOut[21][9][w-1];
              unloadMuxOut[30] = fifoOut[22][9][w-1];
              unloadMuxOut[31] = fifoOut[23][9][w-1];
       end
       16: begin
              unloadMuxOut[0] = fifoOut[24][9][w-1];
              unloadMuxOut[1] = fifoOut[25][9][w-1];
              unloadMuxOut[2] = fifoOut[0][8][w-1];
              unloadMuxOut[3] = fifoOut[1][8][w-1];
              unloadMuxOut[4] = fifoOut[2][8][w-1];
              unloadMuxOut[5] = fifoOut[3][8][w-1];
              unloadMuxOut[6] = fifoOut[4][8][w-1];
              unloadMuxOut[7] = fifoOut[5][8][w-1];
              unloadMuxOut[8] = fifoOut[6][8][w-1];
              unloadMuxOut[9] = fifoOut[7][8][w-1];
              unloadMuxOut[10] = fifoOut[8][8][w-1];
              unloadMuxOut[11] = fifoOut[9][8][w-1];
              unloadMuxOut[12] = fifoOut[10][8][w-1];
              unloadMuxOut[13] = fifoOut[11][8][w-1];
              unloadMuxOut[14] = fifoOut[12][8][w-1];
              unloadMuxOut[15] = fifoOut[13][8][w-1];
              unloadMuxOut[16] = fifoOut[14][8][w-1];
              unloadMuxOut[17] = fifoOut[15][8][w-1];
              unloadMuxOut[18] = fifoOut[16][8][w-1];
              unloadMuxOut[19] = fifoOut[17][8][w-1];
              unloadMuxOut[20] = fifoOut[18][8][w-1];
              unloadMuxOut[21] = fifoOut[19][8][w-1];
              unloadMuxOut[22] = fifoOut[20][8][w-1];
              unloadMuxOut[23] = fifoOut[21][8][w-1];
              unloadMuxOut[24] = fifoOut[22][8][w-1];
              unloadMuxOut[25] = fifoOut[23][8][w-1];
              unloadMuxOut[26] = fifoOut[24][8][w-1];
              unloadMuxOut[27] = fifoOut[25][8][w-1];
              unloadMuxOut[28] = fifoOut[0][7][w-1];
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0;
             end
       end
    endcase
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[38][3];
              muxOutConnector[27] = fifoOut[39][3];
              muxOutConnector[28] = fifoOut[40][3];
              muxOutConnector[29] = fifoOut[41][3];
              muxOutConnector[30] = fifoOut[42][3];
              muxOutConnector[31] = fifoOut[43][3];
              muxOutConnector[32] = fifoOut[44][3];
              muxOutConnector[33] = fifoOut[45][3];
              muxOutConnector[34] = fifoOut[46][3];
              muxOutConnector[35] = fifoOut[47][3];
              muxOutConnector[36] = fifoOut[48][3];
              muxOutConnector[37] = fifoOut[49][3];
              muxOutConnector[38] = fifoOut[50][3];
              muxOutConnector[39] = fifoOut[51][3];
              muxOutConnector[40] = fifoOut[26][2];
              muxOutConnector[41] = fifoOut[27][2];
              muxOutConnector[42] = fifoOut[28][2];
              muxOutConnector[43] = fifoOut[29][2];
              muxOutConnector[44] = fifoOut[30][2];
              muxOutConnector[45] = fifoOut[31][2];
              muxOutConnector[46] = fifoOut[32][2];
              muxOutConnector[47] = fifoOut[33][2];
              muxOutConnector[48] = fifoOut[34][2];
              muxOutConnector[49] = fifoOut[35][2];
              muxOutConnector[50] = fifoOut[36][2];
              muxOutConnector[51] = fifoOut[37][2];
       end
       1: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[38][3];
              muxOutConnector[27] = fifoOut[39][3];
              muxOutConnector[28] = fifoOut[40][3];
              muxOutConnector[29] = fifoOut[41][3];
              muxOutConnector[30] = fifoOut[42][3];
              muxOutConnector[31] = fifoOut[43][3];
              muxOutConnector[32] = fifoOut[44][3];
              muxOutConnector[33] = fifoOut[45][3];
              muxOutConnector[34] = fifoOut[46][3];
              muxOutConnector[35] = fifoOut[47][3];
              muxOutConnector[36] = fifoOut[48][3];
              muxOutConnector[37] = fifoOut[49][3];
              muxOutConnector[38] = fifoOut[50][3];
              muxOutConnector[39] = fifoOut[51][3];
              muxOutConnector[40] = fifoOut[26][2];
              muxOutConnector[41] = fifoOut[27][2];
              muxOutConnector[42] = fifoOut[28][2];
              muxOutConnector[43] = fifoOut[29][2];
              muxOutConnector[44] = fifoOut[30][2];
              muxOutConnector[45] = fifoOut[31][2];
              muxOutConnector[46] = fifoOut[32][2];
              muxOutConnector[47] = fifoOut[33][2];
              muxOutConnector[48] = fifoOut[34][2];
              muxOutConnector[49] = fifoOut[35][2];
              muxOutConnector[50] = fifoOut[36][2];
              muxOutConnector[51] = fifoOut[37][2];
       end
       2: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[38][3];
              muxOutConnector[27] = fifoOut[39][3];
              muxOutConnector[28] = fifoOut[40][3];
              muxOutConnector[29] = fifoOut[41][3];
              muxOutConnector[30] = fifoOut[42][3];
              muxOutConnector[31] = fifoOut[43][3];
              muxOutConnector[32] = fifoOut[44][3];
              muxOutConnector[33] = fifoOut[45][3];
              muxOutConnector[34] = fifoOut[46][3];
              muxOutConnector[35] = fifoOut[47][3];
              muxOutConnector[36] = fifoOut[48][3];
              muxOutConnector[37] = fifoOut[49][3];
              muxOutConnector[38] = fifoOut[50][3];
              muxOutConnector[39] = fifoOut[51][3];
              muxOutConnector[40] = fifoOut[26][2];
              muxOutConnector[41] = fifoOut[27][2];
              muxOutConnector[42] = fifoOut[28][2];
              muxOutConnector[43] = fifoOut[29][2];
              muxOutConnector[44] = fifoOut[30][2];
              muxOutConnector[45] = fifoOut[31][2];
              muxOutConnector[46] = fifoOut[32][2];
              muxOutConnector[47] = fifoOut[33][2];
              muxOutConnector[48] = fifoOut[34][2];
              muxOutConnector[49] = fifoOut[35][2];
              muxOutConnector[50] = fifoOut[36][2];
              muxOutConnector[51] = fifoOut[37][2];
       end
       3: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[38][3];
              muxOutConnector[27] = fifoOut[39][3];
              muxOutConnector[28] = fifoOut[40][3];
              muxOutConnector[29] = fifoOut[41][3];
              muxOutConnector[30] = fifoOut[42][3];
              muxOutConnector[31] = fifoOut[3][2];
              muxOutConnector[32] = fifoOut[4][2];
              muxOutConnector[33] = fifoOut[5][2];
              muxOutConnector[34] = fifoOut[6][2];
              muxOutConnector[35] = fifoOut[7][2];
              muxOutConnector[36] = fifoOut[8][2];
              muxOutConnector[37] = fifoOut[9][2];
              muxOutConnector[38] = fifoOut[10][2];
              muxOutConnector[39] = fifoOut[11][2];
              muxOutConnector[40] = fifoOut[12][2];
              muxOutConnector[41] = fifoOut[13][2];
              muxOutConnector[42] = fifoOut[14][2];
              muxOutConnector[43] = fifoOut[15][2];
              muxOutConnector[44] = fifoOut[16][2];
              muxOutConnector[45] = fifoOut[17][2];
              muxOutConnector[46] = fifoOut[18][2];
              muxOutConnector[47] = fifoOut[19][2];
              muxOutConnector[48] = fifoOut[20][2];
              muxOutConnector[49] = fifoOut[21][2];
              muxOutConnector[50] = fifoOut[22][2];
              muxOutConnector[51] = fifoOut[23][2];
       end
       4: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[24][3];
              muxOutConnector[27] = fifoOut[25][3];
              muxOutConnector[28] = fifoOut[0][2];
              muxOutConnector[29] = fifoOut[1][2];
              muxOutConnector[30] = fifoOut[2][2];
              muxOutConnector[31] = fifoOut[3][2];
              muxOutConnector[32] = fifoOut[4][2];
              muxOutConnector[33] = fifoOut[5][2];
              muxOutConnector[34] = fifoOut[6][2];
              muxOutConnector[35] = fifoOut[7][2];
              muxOutConnector[36] = fifoOut[8][2];
              muxOutConnector[37] = fifoOut[9][2];
              muxOutConnector[38] = fifoOut[10][2];
              muxOutConnector[39] = fifoOut[11][2];
              muxOutConnector[40] = fifoOut[12][2];
              muxOutConnector[41] = fifoOut[13][2];
              muxOutConnector[42] = fifoOut[14][2];
              muxOutConnector[43] = fifoOut[15][2];
              muxOutConnector[44] = fifoOut[16][2];
              muxOutConnector[45] = fifoOut[17][2];
              muxOutConnector[46] = fifoOut[18][2];
              muxOutConnector[47] = fifoOut[19][2];
              muxOutConnector[48] = fifoOut[20][2];
              muxOutConnector[49] = fifoOut[21][2];
              muxOutConnector[50] = fifoOut[22][2];
              muxOutConnector[51] = fifoOut[23][2];
       end
       5: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[24][3];
              muxOutConnector[27] = fifoOut[25][3];
              muxOutConnector[28] = fifoOut[0][2];
              muxOutConnector[29] = fifoOut[1][2];
              muxOutConnector[30] = fifoOut[2][2];
              muxOutConnector[31] = fifoOut[3][2];
              muxOutConnector[32] = fifoOut[4][2];
              muxOutConnector[33] = fifoOut[5][2];
              muxOutConnector[34] = fifoOut[6][2];
              muxOutConnector[35] = fifoOut[7][2];
              muxOutConnector[36] = fifoOut[8][2];
              muxOutConnector[37] = fifoOut[9][2];
              muxOutConnector[38] = fifoOut[10][2];
              muxOutConnector[39] = fifoOut[11][2];
              muxOutConnector[40] = fifoOut[12][2];
              muxOutConnector[41] = fifoOut[13][2];
              muxOutConnector[42] = fifoOut[14][2];
              muxOutConnector[43] = fifoOut[15][2];
              muxOutConnector[44] = fifoOut[16][2];
              muxOutConnector[45] = fifoOut[17][2];
              muxOutConnector[46] = fifoOut[18][2];
              muxOutConnector[47] = fifoOut[19][2];
              muxOutConnector[48] = fifoOut[20][2];
              muxOutConnector[49] = fifoOut[21][2];
              muxOutConnector[50] = fifoOut[22][2];
              muxOutConnector[51] = fifoOut[23][2];
       end
       6: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[17][7];
              muxOutConnector[17] = fifoOut[18][7];
              muxOutConnector[18] = fifoOut[19][7];
              muxOutConnector[19] = fifoOut[20][7];
              muxOutConnector[20] = fifoOut[21][7];
              muxOutConnector[21] = fifoOut[22][7];
              muxOutConnector[22] = fifoOut[23][7];
              muxOutConnector[23] = fifoOut[24][7];
              muxOutConnector[24] = fifoOut[25][7];
              muxOutConnector[25] = fifoOut[0][6];
              muxOutConnector[26] = fifoOut[24][3];
              muxOutConnector[27] = fifoOut[25][3];
              muxOutConnector[28] = fifoOut[0][2];
              muxOutConnector[29] = fifoOut[1][2];
              muxOutConnector[30] = fifoOut[2][2];
              muxOutConnector[31] = fifoOut[3][2];
              muxOutConnector[32] = fifoOut[4][2];
              muxOutConnector[33] = fifoOut[5][2];
              muxOutConnector[34] = fifoOut[6][2];
              muxOutConnector[35] = fifoOut[7][2];
              muxOutConnector[36] = fifoOut[8][2];
              muxOutConnector[37] = fifoOut[9][2];
              muxOutConnector[38] = fifoOut[10][2];
              muxOutConnector[39] = fifoOut[11][2];
              muxOutConnector[40] = fifoOut[12][2];
              muxOutConnector[41] = fifoOut[13][2];
              muxOutConnector[42] = fifoOut[14][2];
              muxOutConnector[43] = fifoOut[15][2];
              muxOutConnector[44] = fifoOut[16][2];
              muxOutConnector[45] = fifoOut[17][2];
              muxOutConnector[46] = fifoOut[18][2];
              muxOutConnector[47] = fifoOut[19][2];
              muxOutConnector[48] = fifoOut[20][2];
              muxOutConnector[49] = fifoOut[21][2];
              muxOutConnector[50] = fifoOut[22][2];
              muxOutConnector[51] = fifoOut[23][2];
       end
       7: begin
              muxOutConnector[0] = fifoOut[1][7];
              muxOutConnector[1] = fifoOut[2][7];
              muxOutConnector[2] = fifoOut[3][7];
              muxOutConnector[3] = fifoOut[4][7];
              muxOutConnector[4] = fifoOut[5][7];
              muxOutConnector[5] = fifoOut[6][7];
              muxOutConnector[6] = fifoOut[7][7];
              muxOutConnector[7] = fifoOut[8][7];
              muxOutConnector[8] = fifoOut[9][7];
              muxOutConnector[9] = fifoOut[10][7];
              muxOutConnector[10] = fifoOut[11][7];
              muxOutConnector[11] = fifoOut[12][7];
              muxOutConnector[12] = fifoOut[13][7];
              muxOutConnector[13] = fifoOut[14][7];
              muxOutConnector[14] = fifoOut[15][7];
              muxOutConnector[15] = fifoOut[16][7];
              muxOutConnector[16] = fifoOut[40][5];
              muxOutConnector[17] = fifoOut[41][5];
              muxOutConnector[18] = fifoOut[42][5];
              muxOutConnector[19] = fifoOut[43][5];
              muxOutConnector[20] = fifoOut[44][5];
              muxOutConnector[21] = fifoOut[45][5];
              muxOutConnector[22] = fifoOut[46][5];
              muxOutConnector[23] = fifoOut[47][5];
              muxOutConnector[24] = fifoOut[48][5];
              muxOutConnector[25] = fifoOut[49][5];
              muxOutConnector[26] = fifoOut[24][3];
              muxOutConnector[27] = fifoOut[25][3];
              muxOutConnector[28] = fifoOut[0][2];
              muxOutConnector[29] = fifoOut[1][2];
              muxOutConnector[30] = fifoOut[2][2];
              muxOutConnector[31] = fifoOut[3][2];
              muxOutConnector[32] = fifoOut[4][2];
              muxOutConnector[33] = fifoOut[5][2];
              muxOutConnector[34] = fifoOut[6][2];
              muxOutConnector[35] = fifoOut[7][2];
              muxOutConnector[36] = fifoOut[8][2];
              muxOutConnector[37] = fifoOut[9][2];
              muxOutConnector[38] = fifoOut[10][2];
              muxOutConnector[39] = fifoOut[11][2];
              muxOutConnector[40] = fifoOut[12][2];
              muxOutConnector[41] = fifoOut[13][2];
              muxOutConnector[42] = fifoOut[14][2];
              muxOutConnector[43] = fifoOut[15][2];
              muxOutConnector[44] = fifoOut[16][2];
              muxOutConnector[45] = fifoOut[17][2];
              muxOutConnector[46] = fifoOut[18][2];
              muxOutConnector[47] = fifoOut[19][2];
              muxOutConnector[48] = fifoOut[20][2];
              muxOutConnector[49] = fifoOut[21][2];
              muxOutConnector[50] = fifoOut[22][2];
              muxOutConnector[51] = fifoOut[23][2];
       end
       8: begin
              muxOutConnector[0] = fifoOut[50][6];
              muxOutConnector[1] = fifoOut[51][6];
              muxOutConnector[2] = fifoOut[26][5];
              muxOutConnector[3] = fifoOut[27][5];
              muxOutConnector[4] = fifoOut[28][5];
              muxOutConnector[5] = fifoOut[29][5];
              muxOutConnector[6] = fifoOut[30][5];
              muxOutConnector[7] = fifoOut[31][5];
              muxOutConnector[8] = fifoOut[32][5];
              muxOutConnector[9] = fifoOut[33][5];
              muxOutConnector[10] = fifoOut[34][5];
              muxOutConnector[11] = fifoOut[35][5];
              muxOutConnector[12] = fifoOut[36][5];
              muxOutConnector[13] = fifoOut[37][5];
              muxOutConnector[14] = fifoOut[38][5];
              muxOutConnector[15] = fifoOut[39][5];
              muxOutConnector[16] = fifoOut[40][5];
              muxOutConnector[17] = fifoOut[41][5];
              muxOutConnector[18] = fifoOut[42][5];
              muxOutConnector[19] = fifoOut[43][5];
              muxOutConnector[20] = fifoOut[44][5];
              muxOutConnector[21] = fifoOut[45][5];
              muxOutConnector[22] = fifoOut[46][5];
              muxOutConnector[23] = fifoOut[47][5];
              muxOutConnector[24] = fifoOut[48][5];
              muxOutConnector[25] = fifoOut[49][5];
              muxOutConnector[26] = fifoOut[24][3];
              muxOutConnector[27] = fifoOut[25][3];
              muxOutConnector[28] = fifoOut[0][2];
              muxOutConnector[29] = fifoOut[1][2];
              muxOutConnector[30] = fifoOut[2][2];
              muxOutConnector[31] = fifoOut[3][2];
              muxOutConnector[32] = fifoOut[4][2];
              muxOutConnector[33] = fifoOut[5][2];
              muxOutConnector[34] = fifoOut[6][2];
              muxOutConnector[35] = fifoOut[7][2];
              muxOutConnector[36] = fifoOut[8][2];
              muxOutConnector[37] = fifoOut[9][2];
              muxOutConnector[38] = fifoOut[10][2];
              muxOutConnector[39] = fifoOut[11][2];
              muxOutConnector[40] = fifoOut[12][2];
              muxOutConnector[41] = fifoOut[13][2];
              muxOutConnector[42] = fifoOut[14][2];
              muxOutConnector[43] = fifoOut[15][2];
              muxOutConnector[44] = fifoOut[16][2];
              muxOutConnector[45] = fifoOut[17][2];
              muxOutConnector[46] = fifoOut[18][2];
              muxOutConnector[47] = fifoOut[19][2];
              muxOutConnector[48] = fifoOut[20][2];
              muxOutConnector[49] = fifoOut[21][2];
              muxOutConnector[50] = fifoOut[22][2];
              muxOutConnector[51] = fifoOut[23][2];
       end
       9: begin
              muxOutConnector[0] = fifoOut[50][6];
              muxOutConnector[1] = fifoOut[51][6];
              muxOutConnector[2] = fifoOut[26][5];
              muxOutConnector[3] = fifoOut[27][5];
              muxOutConnector[4] = fifoOut[28][5];
              muxOutConnector[5] = fifoOut[29][5];
              muxOutConnector[6] = fifoOut[30][5];
              muxOutConnector[7] = fifoOut[31][5];
              muxOutConnector[8] = fifoOut[32][5];
              muxOutConnector[9] = fifoOut[33][5];
              muxOutConnector[10] = fifoOut[34][5];
              muxOutConnector[11] = fifoOut[35][5];
              muxOutConnector[12] = fifoOut[36][5];
              muxOutConnector[13] = fifoOut[37][5];
              muxOutConnector[14] = fifoOut[38][5];
              muxOutConnector[15] = fifoOut[39][5];
              muxOutConnector[16] = fifoOut[40][5];
              muxOutConnector[17] = fifoOut[41][5];
              muxOutConnector[18] = fifoOut[42][5];
              muxOutConnector[19] = fifoOut[43][5];
              muxOutConnector[20] = fifoOut[44][5];
              muxOutConnector[21] = fifoOut[45][5];
              muxOutConnector[22] = fifoOut[46][5];
              muxOutConnector[23] = fifoOut[47][5];
              muxOutConnector[24] = fifoOut[48][5];
              muxOutConnector[25] = fifoOut[49][5];
              muxOutConnector[26] = fifoOut[24][3];
              muxOutConnector[27] = fifoOut[25][3];
              muxOutConnector[28] = fifoOut[0][2];
              muxOutConnector[29] = fifoOut[1][2];
              muxOutConnector[30] = fifoOut[2][2];
              muxOutConnector[31] = fifoOut[3][2];
              muxOutConnector[32] = fifoOut[4][2];
              muxOutConnector[33] = fifoOut[5][2];
              muxOutConnector[34] = fifoOut[6][2];
              muxOutConnector[35] = fifoOut[7][2];
              muxOutConnector[36] = fifoOut[8][2];
              muxOutConnector[37] = fifoOut[9][2];
              muxOutConnector[38] = fifoOut[10][2];
              muxOutConnector[39] = fifoOut[11][2];
              muxOutConnector[40] = fifoOut[12][2];
              muxOutConnector[41] = fifoOut[13][2];
              muxOutConnector[42] = fifoOut[14][2];
              muxOutConnector[43] = fifoOut[15][2];
              muxOutConnector[44] = fifoOut[16][2];
              muxOutConnector[45] = fifoOut[17][2];
              muxOutConnector[46] = fifoOut[18][2];
              muxOutConnector[47] = fifoOut[19][2];
              muxOutConnector[48] = fifoOut[20][2];
              muxOutConnector[49] = fifoOut[21][2];
              muxOutConnector[50] = fifoOut[22][2];
              muxOutConnector[51] = fifoOut[23][2];
       end
       10: begin
              muxOutConnector[0] = fifoOut[50][6];
              muxOutConnector[1] = fifoOut[51][6];
              muxOutConnector[2] = fifoOut[26][5];
              muxOutConnector[3] = fifoOut[27][5];
              muxOutConnector[4] = fifoOut[28][5];
              muxOutConnector[5] = fifoOut[29][5];
              muxOutConnector[6] = fifoOut[30][5];
              muxOutConnector[7] = fifoOut[31][5];
              muxOutConnector[8] = fifoOut[32][5];
              muxOutConnector[9] = fifoOut[33][5];
              muxOutConnector[10] = fifoOut[34][5];
              muxOutConnector[11] = fifoOut[35][5];
              muxOutConnector[12] = fifoOut[36][5];
              muxOutConnector[13] = fifoOut[37][5];
              muxOutConnector[14] = fifoOut[38][5];
              muxOutConnector[15] = fifoOut[39][5];
              muxOutConnector[16] = fifoOut[40][5];
              muxOutConnector[17] = fifoOut[41][5];
              muxOutConnector[18] = fifoOut[42][5];
              muxOutConnector[19] = fifoOut[43][5];
              muxOutConnector[20] = fifoOut[44][5];
              muxOutConnector[21] = fifoOut[45][5];
              muxOutConnector[22] = fifoOut[46][5];
              muxOutConnector[23] = fifoOut[47][5];
              muxOutConnector[24] = fifoOut[48][5];
              muxOutConnector[25] = fifoOut[49][5];
              muxOutConnector[26] = fifoOut[24][3];
              muxOutConnector[27] = fifoOut[25][3];
              muxOutConnector[28] = fifoOut[0][2];
              muxOutConnector[29] = fifoOut[1][2];
              muxOutConnector[30] = fifoOut[2][2];
              muxOutConnector[31] = fifoOut[3][2];
              muxOutConnector[32] = fifoOut[4][2];
              muxOutConnector[33] = fifoOut[5][2];
              muxOutConnector[34] = fifoOut[6][2];
              muxOutConnector[35] = fifoOut[7][2];
              muxOutConnector[36] = fifoOut[8][2];
              muxOutConnector[37] = fifoOut[9][2];
              muxOutConnector[38] = fifoOut[10][2];
              muxOutConnector[39] = fifoOut[11][2];
              muxOutConnector[40] = fifoOut[12][2];
              muxOutConnector[41] = fifoOut[13][2];
              muxOutConnector[42] = fifoOut[14][2];
              muxOutConnector[43] = fifoOut[15][2];
              muxOutConnector[44] = fifoOut[16][2];
              muxOutConnector[45] = fifoOut[17][2];
              muxOutConnector[46] = fifoOut[18][2];
              muxOutConnector[47] = fifoOut[19][2];
              muxOutConnector[48] = fifoOut[20][2];
              muxOutConnector[49] = fifoOut[21][2];
              muxOutConnector[50] = fifoOut[22][2];
              muxOutConnector[51] = fifoOut[23][2];
       end
       11: begin
              muxOutConnector[0] = fifoOut[50][6];
              muxOutConnector[1] = fifoOut[51][6];
              muxOutConnector[2] = fifoOut[26][5];
              muxOutConnector[3] = fifoOut[27][5];
              muxOutConnector[4] = fifoOut[28][5];
              muxOutConnector[5] = fifoOut[29][5];
              muxOutConnector[6] = fifoOut[30][5];
              muxOutConnector[7] = fifoOut[31][5];
              muxOutConnector[8] = fifoOut[32][5];
              muxOutConnector[9] = fifoOut[33][5];
              muxOutConnector[10] = fifoOut[34][5];
              muxOutConnector[11] = fifoOut[35][5];
              muxOutConnector[12] = fifoOut[36][5];
              muxOutConnector[13] = fifoOut[37][5];
              muxOutConnector[14] = fifoOut[38][5];
              muxOutConnector[15] = fifoOut[39][5];
              muxOutConnector[16] = fifoOut[40][5];
              muxOutConnector[17] = fifoOut[41][5];
              muxOutConnector[18] = fifoOut[42][5];
              muxOutConnector[19] = fifoOut[43][5];
              muxOutConnector[20] = fifoOut[44][5];
              muxOutConnector[21] = fifoOut[45][5];
              muxOutConnector[22] = fifoOut[46][5];
              muxOutConnector[23] = fifoOut[47][5];
              muxOutConnector[24] = fifoOut[48][5];
              muxOutConnector[25] = fifoOut[49][5];
              muxOutConnector[26] = fifoOut[24][3];
              muxOutConnector[27] = fifoOut[25][3];
              muxOutConnector[28] = fifoOut[0][2];
              muxOutConnector[29] = fifoOut[1][2];
              muxOutConnector[30] = fifoOut[2][2];
              muxOutConnector[31] = fifoOut[3][2];
              muxOutConnector[32] = fifoOut[4][2];
              muxOutConnector[33] = fifoOut[5][2];
              muxOutConnector[34] = fifoOut[6][2];
              muxOutConnector[35] = fifoOut[7][2];
              muxOutConnector[36] = fifoOut[8][2];
              muxOutConnector[37] = fifoOut[9][2];
              muxOutConnector[38] = fifoOut[10][2];
              muxOutConnector[39] = fifoOut[11][2];
              muxOutConnector[40] = fifoOut[12][2];
              muxOutConnector[41] = fifoOut[13][2];
              muxOutConnector[42] = fifoOut[14][2];
              muxOutConnector[43] = fifoOut[15][2];
              muxOutConnector[44] = fifoOut[16][2];
              muxOutConnector[45] = fifoOut[17][2];
              muxOutConnector[46] = fifoOut[18][2];
              muxOutConnector[47] = fifoOut[19][2];
              muxOutConnector[48] = fifoOut[20][2];
              muxOutConnector[49] = fifoOut[21][2];
              muxOutConnector[50] = fifoOut[22][2];
              muxOutConnector[51] = fifoOut[23][2];
       end
       12: begin
              muxOutConnector[0] = fifoOut[50][6];
              muxOutConnector[1] = fifoOut[51][6];
              muxOutConnector[2] = fifoOut[26][5];
              muxOutConnector[3] = fifoOut[27][5];
              muxOutConnector[4] = fifoOut[28][5];
              muxOutConnector[5] = fifoOut[29][5];
              muxOutConnector[6] = fifoOut[30][5];
              muxOutConnector[7] = fifoOut[31][5];
              muxOutConnector[8] = fifoOut[32][5];
              muxOutConnector[9] = fifoOut[33][5];
              muxOutConnector[10] = fifoOut[34][5];
              muxOutConnector[11] = fifoOut[35][5];
              muxOutConnector[12] = fifoOut[36][5];
              muxOutConnector[13] = fifoOut[37][5];
              muxOutConnector[14] = fifoOut[38][5];
              muxOutConnector[15] = fifoOut[39][5];
              muxOutConnector[16] = fifoOut[40][5];
              muxOutConnector[17] = fifoOut[41][5];
              muxOutConnector[18] = fifoOut[42][5];
              muxOutConnector[19] = fifoOut[43][5];
              muxOutConnector[20] = fifoOut[44][5];
              muxOutConnector[21] = fifoOut[45][5];
              muxOutConnector[22] = fifoOut[46][5];
              muxOutConnector[23] = fifoOut[47][5];
              muxOutConnector[24] = fifoOut[48][5];
              muxOutConnector[25] = fifoOut[49][5];
              muxOutConnector[26] = fifoOut[24][3];
              muxOutConnector[27] = fifoOut[25][3];
              muxOutConnector[28] = fifoOut[0][2];
              muxOutConnector[29] = fifoOut[1][2];
              muxOutConnector[30] = fifoOut[2][2];
              muxOutConnector[31] = fifoOut[3][2];
              muxOutConnector[32] = fifoOut[4][2];
              muxOutConnector[33] = fifoOut[5][2];
              muxOutConnector[34] = fifoOut[6][2];
              muxOutConnector[35] = fifoOut[7][2];
              muxOutConnector[36] = fifoOut[8][2];
              muxOutConnector[37] = fifoOut[9][2];
              muxOutConnector[38] = fifoOut[10][2];
              muxOutConnector[39] = fifoOut[11][2];
              muxOutConnector[40] = fifoOut[12][2];
              muxOutConnector[41] = fifoOut[13][2];
              muxOutConnector[42] = fifoOut[14][2];
              muxOutConnector[43] = fifoOut[15][2];
              muxOutConnector[44] = fifoOut[16][2];
              muxOutConnector[45] = fifoOut[17][2];
              muxOutConnector[46] = fifoOut[18][2];
              muxOutConnector[47] = fifoOut[19][2];
              muxOutConnector[48] = fifoOut[20][2];
              muxOutConnector[49] = fifoOut[21][2];
              muxOutConnector[50] = fifoOut[22][2];
              muxOutConnector[51] = fifoOut[23][2];
       end
       13: begin
              muxOutConnector[0] = fifoOut[50][6];
              muxOutConnector[1] = fifoOut[51][6];
              muxOutConnector[2] = fifoOut[26][5];
              muxOutConnector[3] = fifoOut[27][5];
              muxOutConnector[4] = fifoOut[28][5];
              muxOutConnector[5] = fifoOut[29][5];
              muxOutConnector[6] = fifoOut[30][5];
              muxOutConnector[7] = fifoOut[31][5];
              muxOutConnector[8] = fifoOut[32][5];
              muxOutConnector[9] = fifoOut[33][5];
              muxOutConnector[10] = fifoOut[34][5];
              muxOutConnector[11] = fifoOut[35][5];
              muxOutConnector[12] = fifoOut[36][5];
              muxOutConnector[13] = fifoOut[37][5];
              muxOutConnector[14] = fifoOut[38][5];
              muxOutConnector[15] = fifoOut[39][5];
              muxOutConnector[16] = fifoOut[40][5];
              muxOutConnector[17] = fifoOut[41][5];
              muxOutConnector[18] = fifoOut[42][5];
              muxOutConnector[19] = fifoOut[43][5];
              muxOutConnector[20] = fifoOut[44][5];
              muxOutConnector[21] = fifoOut[45][5];
              muxOutConnector[22] = fifoOut[46][5];
              muxOutConnector[23] = fifoOut[47][5];
              muxOutConnector[24] = fifoOut[48][5];
              muxOutConnector[25] = fifoOut[49][5];
              muxOutConnector[26] = fifoOut[24][3];
              muxOutConnector[27] = fifoOut[25][3];
              muxOutConnector[28] = fifoOut[0][2];
              muxOutConnector[29] = fifoOut[1][2];
              muxOutConnector[30] = fifoOut[2][2];
              muxOutConnector[31] = fifoOut[3][2];
              muxOutConnector[32] = fifoOut[4][2];
              muxOutConnector[33] = fifoOut[5][2];
              muxOutConnector[34] = fifoOut[6][2];
              muxOutConnector[35] = fifoOut[7][2];
              muxOutConnector[36] = fifoOut[8][2];
              muxOutConnector[37] = fifoOut[9][2];
              muxOutConnector[38] = fifoOut[10][2];
              muxOutConnector[39] = fifoOut[11][2];
              muxOutConnector[40] = fifoOut[12][2];
              muxOutConnector[41] = fifoOut[13][2];
              muxOutConnector[42] = fifoOut[14][2];
              muxOutConnector[43] = fifoOut[15][2];
              muxOutConnector[44] = fifoOut[16][2];
              muxOutConnector[45] = fifoOut[40][0];
              muxOutConnector[46] = fifoOut[41][0];
              muxOutConnector[47] = fifoOut[42][0];
              muxOutConnector[48] = fifoOut[43][0];
              muxOutConnector[49] = fifoOut[44][0];
              muxOutConnector[50] = fifoOut[45][0];
              muxOutConnector[51] = fifoOut[46][0];
       end
       14: begin
              muxOutConnector[0] = fifoOut[50][6];
              muxOutConnector[1] = fifoOut[51][6];
              muxOutConnector[2] = fifoOut[26][5];
              muxOutConnector[3] = fifoOut[27][5];
              muxOutConnector[4] = fifoOut[28][5];
              muxOutConnector[5] = fifoOut[29][5];
              muxOutConnector[6] = fifoOut[30][5];
              muxOutConnector[7] = fifoOut[31][5];
              muxOutConnector[8] = fifoOut[32][5];
              muxOutConnector[9] = fifoOut[33][5];
              muxOutConnector[10] = fifoOut[34][5];
              muxOutConnector[11] = fifoOut[35][5];
              muxOutConnector[12] = fifoOut[36][5];
              muxOutConnector[13] = fifoOut[37][5];
              muxOutConnector[14] = fifoOut[38][5];
              muxOutConnector[15] = fifoOut[39][5];
              muxOutConnector[16] = fifoOut[40][5];
              muxOutConnector[17] = fifoOut[41][5];
              muxOutConnector[18] = fifoOut[42][5];
              muxOutConnector[19] = fifoOut[43][5];
              muxOutConnector[20] = fifoOut[44][5];
              muxOutConnector[21] = fifoOut[45][5];
              muxOutConnector[22] = fifoOut[46][5];
              muxOutConnector[23] = fifoOut[47][5];
              muxOutConnector[24] = fifoOut[48][5];
              muxOutConnector[25] = fifoOut[49][5];
              muxOutConnector[26] = fifoOut[47][1];
              muxOutConnector[27] = fifoOut[48][1];
              muxOutConnector[28] = fifoOut[49][1];
              muxOutConnector[29] = fifoOut[50][1];
              muxOutConnector[30] = fifoOut[51][1];
              muxOutConnector[31] = fifoOut[26][0];
              muxOutConnector[32] = fifoOut[27][0];
              muxOutConnector[33] = fifoOut[28][0];
              muxOutConnector[34] = fifoOut[29][0];
              muxOutConnector[35] = fifoOut[30][0];
              muxOutConnector[36] = fifoOut[31][0];
              muxOutConnector[37] = fifoOut[32][0];
              muxOutConnector[38] = fifoOut[33][0];
              muxOutConnector[39] = fifoOut[34][0];
              muxOutConnector[40] = fifoOut[35][0];
              muxOutConnector[41] = fifoOut[36][0];
              muxOutConnector[42] = fifoOut[37][0];
              muxOutConnector[43] = fifoOut[38][0];
              muxOutConnector[44] = fifoOut[39][0];
              muxOutConnector[45] = fifoOut[40][0];
              muxOutConnector[46] = fifoOut[41][0];
              muxOutConnector[47] = fifoOut[42][0];
              muxOutConnector[48] = fifoOut[43][0];
              muxOutConnector[49] = fifoOut[44][0];
              muxOutConnector[50] = fifoOut[45][0];
              muxOutConnector[51] = fifoOut[46][0];
       end
       15: begin
              muxOutConnector[0] = fifoOut[50][6];
              muxOutConnector[1] = fifoOut[51][6];
              muxOutConnector[2] = fifoOut[26][5];
              muxOutConnector[3] = fifoOut[27][5];
              muxOutConnector[4] = fifoOut[28][5];
              muxOutConnector[5] = fifoOut[29][5];
              muxOutConnector[6] = fifoOut[30][5];
              muxOutConnector[7] = fifoOut[31][5];
              muxOutConnector[8] = fifoOut[32][5];
              muxOutConnector[9] = fifoOut[33][5];
              muxOutConnector[10] = fifoOut[34][5];
              muxOutConnector[11] = fifoOut[35][5];
              muxOutConnector[12] = fifoOut[36][5];
              muxOutConnector[13] = fifoOut[37][5];
              muxOutConnector[14] = fifoOut[38][5];
              muxOutConnector[15] = fifoOut[39][5];
              muxOutConnector[16] = fifoOut[40][5];
              muxOutConnector[17] = fifoOut[41][5];
              muxOutConnector[18] = fifoOut[42][5];
              muxOutConnector[19] = fifoOut[43][5];
              muxOutConnector[20] = fifoOut[44][5];
              muxOutConnector[21] = fifoOut[45][5];
              muxOutConnector[22] = fifoOut[46][5];
              muxOutConnector[23] = fifoOut[47][5];
              muxOutConnector[24] = fifoOut[48][5];
              muxOutConnector[25] = fifoOut[49][5];
              muxOutConnector[26] = fifoOut[47][1];
              muxOutConnector[27] = fifoOut[48][1];
              muxOutConnector[28] = fifoOut[49][1];
              muxOutConnector[29] = fifoOut[50][1];
              muxOutConnector[30] = fifoOut[51][1];
              muxOutConnector[31] = fifoOut[26][0];
              muxOutConnector[32] = fifoOut[27][0];
              muxOutConnector[33] = fifoOut[28][0];
              muxOutConnector[34] = fifoOut[29][0];
              muxOutConnector[35] = fifoOut[30][0];
              muxOutConnector[36] = fifoOut[31][0];
              muxOutConnector[37] = fifoOut[32][0];
              muxOutConnector[38] = fifoOut[33][0];
              muxOutConnector[39] = fifoOut[34][0];
              muxOutConnector[40] = fifoOut[35][0];
              muxOutConnector[41] = fifoOut[36][0];
              muxOutConnector[42] = fifoOut[37][0];
              muxOutConnector[43] = fifoOut[38][0];
              muxOutConnector[44] = fifoOut[39][0];
              muxOutConnector[45] = fifoOut[40][0];
              muxOutConnector[46] = fifoOut[41][0];
              muxOutConnector[47] = fifoOut[42][0];
              muxOutConnector[48] = fifoOut[43][0];
              muxOutConnector[49] = fifoOut[44][0];
              muxOutConnector[50] = fifoOut[45][0];
              muxOutConnector[51] = fifoOut[46][0];
       end
       16: begin
              muxOutConnector[0] = fifoOut[50][6];
              muxOutConnector[1] = fifoOut[51][6];
              muxOutConnector[2] = fifoOut[26][5];
              muxOutConnector[3] = fifoOut[27][5];
              muxOutConnector[4] = fifoOut[28][5];
              muxOutConnector[5] = fifoOut[29][5];
              muxOutConnector[6] = fifoOut[30][5];
              muxOutConnector[7] = fifoOut[31][5];
              muxOutConnector[8] = fifoOut[32][5];
              muxOutConnector[9] = fifoOut[33][5];
              muxOutConnector[10] = fifoOut[34][5];
              muxOutConnector[11] = fifoOut[35][5];
              muxOutConnector[12] = fifoOut[36][5];
              muxOutConnector[13] = fifoOut[37][5];
              muxOutConnector[14] = fifoOut[38][5];
              muxOutConnector[15] = fifoOut[39][5];
              muxOutConnector[16] = fifoOut[40][5];
              muxOutConnector[17] = fifoOut[41][5];
              muxOutConnector[18] = fifoOut[42][5];
              muxOutConnector[19] = fifoOut[3][4];
              muxOutConnector[20] = fifoOut[4][4];
              muxOutConnector[21] = fifoOut[5][4];
              muxOutConnector[22] = fifoOut[6][4];
              muxOutConnector[23] = fifoOut[7][4];
              muxOutConnector[24] = fifoOut[8][4];
              muxOutConnector[25] = fifoOut[9][4];
              muxOutConnector[26] = fifoOut[47][1];
              muxOutConnector[27] = fifoOut[48][1];
              muxOutConnector[28] = fifoOut[49][1];
              muxOutConnector[29] = fifoOut[50][1];
              muxOutConnector[30] = fifoOut[51][1];
              muxOutConnector[31] = fifoOut[26][0];
              muxOutConnector[32] = fifoOut[27][0];
              muxOutConnector[33] = fifoOut[28][0];
              muxOutConnector[34] = fifoOut[29][0];
              muxOutConnector[35] = fifoOut[30][0];
              muxOutConnector[36] = fifoOut[31][0];
              muxOutConnector[37] = fifoOut[32][0];
              muxOutConnector[38] = fifoOut[33][0];
              muxOutConnector[39] = fifoOut[34][0];
              muxOutConnector[40] = fifoOut[35][0];
              muxOutConnector[41] = fifoOut[36][0];
              muxOutConnector[42] = fifoOut[37][0];
              muxOutConnector[43] = fifoOut[38][0];
              muxOutConnector[44] = fifoOut[39][0];
              muxOutConnector[45] = fifoOut[40][0];
              muxOutConnector[46] = fifoOut[41][0];
              muxOutConnector[47] = fifoOut[42][0];
              muxOutConnector[48] = fifoOut[43][0];
              muxOutConnector[49] = fifoOut[44][0];
              muxOutConnector[50] = fifoOut[45][0];
              muxOutConnector[51] = fifoOut[46][0];
       end
       17: begin
              muxOutConnector[0] = fifoOut[10][5];
              muxOutConnector[1] = fifoOut[11][5];
              muxOutConnector[2] = fifoOut[12][5];
              muxOutConnector[3] = fifoOut[13][5];
              muxOutConnector[4] = fifoOut[14][5];
              muxOutConnector[5] = fifoOut[15][5];
              muxOutConnector[6] = fifoOut[16][5];
              muxOutConnector[7] = fifoOut[17][5];
              muxOutConnector[8] = fifoOut[18][5];
              muxOutConnector[9] = fifoOut[19][5];
              muxOutConnector[10] = fifoOut[20][5];
              muxOutConnector[11] = fifoOut[21][5];
              muxOutConnector[12] = fifoOut[22][5];
              muxOutConnector[13] = fifoOut[23][5];
              muxOutConnector[14] = fifoOut[24][5];
              muxOutConnector[15] = fifoOut[25][5];
              muxOutConnector[16] = fifoOut[0][4];
              muxOutConnector[17] = fifoOut[1][4];
              muxOutConnector[18] = fifoOut[2][4];
              muxOutConnector[19] = fifoOut[3][4];
              muxOutConnector[20] = fifoOut[4][4];
              muxOutConnector[21] = fifoOut[5][4];
              muxOutConnector[22] = fifoOut[6][4];
              muxOutConnector[23] = fifoOut[7][4];
              muxOutConnector[24] = fifoOut[8][4];
              muxOutConnector[25] = fifoOut[9][4];
              muxOutConnector[26] = fifoOut[47][1];
              muxOutConnector[27] = fifoOut[48][1];
              muxOutConnector[28] = fifoOut[49][1];
              muxOutConnector[29] = fifoOut[50][1];
              muxOutConnector[30] = fifoOut[51][1];
              muxOutConnector[31] = fifoOut[26][0];
              muxOutConnector[32] = fifoOut[27][0];
              muxOutConnector[33] = fifoOut[28][0];
              muxOutConnector[34] = fifoOut[29][0];
              muxOutConnector[35] = fifoOut[30][0];
              muxOutConnector[36] = fifoOut[31][0];
              muxOutConnector[37] = fifoOut[32][0];
              muxOutConnector[38] = fifoOut[33][0];
              muxOutConnector[39] = fifoOut[34][0];
              muxOutConnector[40] = fifoOut[35][0];
              muxOutConnector[41] = fifoOut[36][0];
              muxOutConnector[42] = fifoOut[37][0];
              muxOutConnector[43] = fifoOut[38][0];
              muxOutConnector[44] = fifoOut[39][0];
              muxOutConnector[45] = fifoOut[40][0];
              muxOutConnector[46] = fifoOut[41][0];
              muxOutConnector[47] = fifoOut[42][0];
              muxOutConnector[48] = fifoOut[43][0];
              muxOutConnector[49] = fifoOut[44][0];
              muxOutConnector[50] = fifoOut[45][0];
              muxOutConnector[51] = fifoOut[46][0];
       end
       18: begin
              muxOutConnector[0] = fifoOut[10][5];
              muxOutConnector[1] = fifoOut[11][5];
              muxOutConnector[2] = fifoOut[12][5];
              muxOutConnector[3] = fifoOut[13][5];
              muxOutConnector[4] = fifoOut[14][5];
              muxOutConnector[5] = fifoOut[15][5];
              muxOutConnector[6] = fifoOut[16][5];
              muxOutConnector[7] = fifoOut[17][5];
              muxOutConnector[8] = fifoOut[18][5];
              muxOutConnector[9] = fifoOut[19][5];
              muxOutConnector[10] = fifoOut[20][5];
              muxOutConnector[11] = fifoOut[21][5];
              muxOutConnector[12] = fifoOut[22][5];
              muxOutConnector[13] = fifoOut[23][5];
              muxOutConnector[14] = fifoOut[24][5];
              muxOutConnector[15] = fifoOut[25][5];
              muxOutConnector[16] = fifoOut[0][4];
              muxOutConnector[17] = fifoOut[1][4];
              muxOutConnector[18] = fifoOut[2][4];
              muxOutConnector[19] = fifoOut[3][4];
              muxOutConnector[20] = fifoOut[4][4];
              muxOutConnector[21] = fifoOut[5][4];
              muxOutConnector[22] = fifoOut[6][4];
              muxOutConnector[23] = fifoOut[7][4];
              muxOutConnector[24] = fifoOut[8][4];
              muxOutConnector[25] = fifoOut[9][4];
              muxOutConnector[26] = fifoOut[47][1];
              muxOutConnector[27] = fifoOut[48][1];
              muxOutConnector[28] = fifoOut[49][1];
              muxOutConnector[29] = fifoOut[50][1];
              muxOutConnector[30] = fifoOut[51][1];
              muxOutConnector[31] = fifoOut[26][0];
              muxOutConnector[32] = fifoOut[27][0];
              muxOutConnector[33] = fifoOut[28][0];
              muxOutConnector[34] = fifoOut[29][0];
              muxOutConnector[35] = fifoOut[30][0];
              muxOutConnector[36] = fifoOut[31][0];
              muxOutConnector[37] = fifoOut[32][0];
              muxOutConnector[38] = fifoOut[33][0];
              muxOutConnector[39] = fifoOut[34][0];
              muxOutConnector[40] = fifoOut[35][0];
              muxOutConnector[41] = fifoOut[36][0];
              muxOutConnector[42] = fifoOut[37][0];
              muxOutConnector[43] = fifoOut[38][0];
              muxOutConnector[44] = fifoOut[39][0];
              muxOutConnector[45] = fifoOut[40][0];
              muxOutConnector[46] = fifoOut[41][0];
              muxOutConnector[47] = fifoOut[42][0];
              muxOutConnector[48] = fifoOut[43][0];
              muxOutConnector[49] = fifoOut[44][0];
              muxOutConnector[50] = fifoOut[45][0];
              muxOutConnector[51] = fifoOut[46][0];
       end
       19: begin
              muxOutConnector[0] = fifoOut[10][5];
              muxOutConnector[1] = fifoOut[11][5];
              muxOutConnector[2] = fifoOut[12][5];
              muxOutConnector[3] = fifoOut[13][5];
              muxOutConnector[4] = fifoOut[14][5];
              muxOutConnector[5] = fifoOut[15][5];
              muxOutConnector[6] = fifoOut[16][5];
              muxOutConnector[7] = fifoOut[17][5];
              muxOutConnector[8] = fifoOut[18][5];
              muxOutConnector[9] = fifoOut[19][5];
              muxOutConnector[10] = fifoOut[20][5];
              muxOutConnector[11] = fifoOut[21][5];
              muxOutConnector[12] = fifoOut[22][5];
              muxOutConnector[13] = fifoOut[23][5];
              muxOutConnector[14] = fifoOut[24][5];
              muxOutConnector[15] = fifoOut[25][5];
              muxOutConnector[16] = fifoOut[0][4];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[47][1];
              muxOutConnector[27] = fifoOut[48][1];
              muxOutConnector[28] = fifoOut[49][1];
              muxOutConnector[29] = fifoOut[50][1];
              muxOutConnector[30] = fifoOut[51][1];
              muxOutConnector[31] = fifoOut[26][0];
              muxOutConnector[32] = fifoOut[27][0];
              muxOutConnector[33] = fifoOut[28][0];
              muxOutConnector[34] = fifoOut[29][0];
              muxOutConnector[35] = fifoOut[30][0];
              muxOutConnector[36] = fifoOut[31][0];
              muxOutConnector[37] = fifoOut[32][0];
              muxOutConnector[38] = fifoOut[33][0];
              muxOutConnector[39] = fifoOut[34][0];
              muxOutConnector[40] = fifoOut[35][0];
              muxOutConnector[41] = fifoOut[36][0];
              muxOutConnector[42] = fifoOut[37][0];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
