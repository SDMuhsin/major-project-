`timescale 1ns / 1ps
module LMem0To1_511_circ0_ys_scripted(
        muxOut,
        ly0In,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 14;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

reg   feedback_en;
reg [ w - 1 : 0 ]column_1[ r - 1 : 0 ];
reg chip_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(chip_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= column_1[i];
         end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
  feedback_en=rd_en;
      if(wr_en)begin
        chip_en=wr_en;
      end
      else begin
        chip_en=feedback_en;
      end
   if(feedback_en)begin
      for(i = r-1; i > -1; i=i-1) begin
        column_1[i] <= fifoOut[i][c-1];
      end
   end
   else begin
      for(i = r-1; i > -1; i=i-1) begin
        column_1[i] <= ly0InConnector[i];
      end
    end
end
always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[44][3];
              muxOutConnector[1] = fifoOut[45][3];
              muxOutConnector[2] = fifoOut[46][3];
              muxOutConnector[3] = fifoOut[47][3];
              muxOutConnector[4] = fifoOut[48][3];
              muxOutConnector[5] = fifoOut[49][3];
              muxOutConnector[6] = fifoOut[50][3];
              muxOutConnector[7] = fifoOut[51][3];
              muxOutConnector[8] = fifoOut[26][2];
              muxOutConnector[9] = fifoOut[27][2];
              muxOutConnector[10] = fifoOut[28][2];
              muxOutConnector[11] = fifoOut[29][2];
              muxOutConnector[12] = fifoOut[30][2];
              muxOutConnector[13] = fifoOut[31][2];
              muxOutConnector[14] = fifoOut[32][2];
              muxOutConnector[15] = fifoOut[33][2];
              muxOutConnector[16] = fifoOut[34][2];
              muxOutConnector[17] = fifoOut[35][2];
              muxOutConnector[18] = fifoOut[36][2];
              muxOutConnector[19] = fifoOut[37][2];
              muxOutConnector[20] = fifoOut[38][2];
              muxOutConnector[21] = fifoOut[39][2];
              muxOutConnector[22] = fifoOut[40][2];
              muxOutConnector[23] = fifoOut[41][2];
              muxOutConnector[24] = fifoOut[42][2];
              muxOutConnector[25] = fifoOut[43][2];
              muxOutConnector[26] = fifoOut[35][8];
              muxOutConnector[27] = fifoOut[36][8];
              muxOutConnector[28] = fifoOut[37][8];
              muxOutConnector[29] = fifoOut[38][8];
              muxOutConnector[30] = fifoOut[39][8];
              muxOutConnector[31] = fifoOut[40][8];
              muxOutConnector[32] = fifoOut[41][8];
              muxOutConnector[33] = fifoOut[42][8];
              muxOutConnector[34] = fifoOut[43][8];
              muxOutConnector[35] = fifoOut[44][8];
              muxOutConnector[36] = fifoOut[45][8];
              muxOutConnector[37] = fifoOut[46][8];
              muxOutConnector[38] = fifoOut[47][8];
              muxOutConnector[39] = fifoOut[48][8];
              muxOutConnector[40] = fifoOut[49][8];
              muxOutConnector[41] = fifoOut[50][8];
              muxOutConnector[42] = fifoOut[51][8];
              muxOutConnector[43] = fifoOut[26][7];
              muxOutConnector[44] = fifoOut[27][7];
              muxOutConnector[45] = fifoOut[28][7];
              muxOutConnector[46] = fifoOut[29][7];
              muxOutConnector[47] = fifoOut[30][7];
              muxOutConnector[48] = fifoOut[31][7];
              muxOutConnector[49] = fifoOut[32][7];
              muxOutConnector[50] = fifoOut[33][7];
              muxOutConnector[51] = fifoOut[34][7];
       end
       1: begin
              muxOutConnector[0] = fifoOut[44][3];
              muxOutConnector[1] = fifoOut[45][3];
              muxOutConnector[2] = fifoOut[46][3];
              muxOutConnector[3] = fifoOut[47][3];
              muxOutConnector[4] = fifoOut[48][3];
              muxOutConnector[5] = fifoOut[49][3];
              muxOutConnector[6] = fifoOut[50][3];
              muxOutConnector[7] = fifoOut[51][3];
              muxOutConnector[8] = fifoOut[26][2];
              muxOutConnector[9] = fifoOut[27][2];
              muxOutConnector[10] = fifoOut[28][2];
              muxOutConnector[11] = fifoOut[29][2];
              muxOutConnector[12] = fifoOut[30][2];
              muxOutConnector[13] = fifoOut[31][2];
              muxOutConnector[14] = fifoOut[32][2];
              muxOutConnector[15] = fifoOut[33][2];
              muxOutConnector[16] = fifoOut[34][2];
              muxOutConnector[17] = fifoOut[35][2];
              muxOutConnector[18] = fifoOut[36][2];
              muxOutConnector[19] = fifoOut[37][2];
              muxOutConnector[20] = fifoOut[38][2];
              muxOutConnector[21] = fifoOut[39][2];
              muxOutConnector[22] = fifoOut[40][2];
              muxOutConnector[23] = fifoOut[41][2];
              muxOutConnector[24] = fifoOut[42][2];
              muxOutConnector[25] = fifoOut[43][2];
              muxOutConnector[26] = fifoOut[35][8];
              muxOutConnector[27] = fifoOut[36][8];
              muxOutConnector[28] = fifoOut[37][8];
              muxOutConnector[29] = fifoOut[38][8];
              muxOutConnector[30] = fifoOut[39][8];
              muxOutConnector[31] = fifoOut[40][8];
              muxOutConnector[32] = fifoOut[41][8];
              muxOutConnector[33] = fifoOut[42][8];
              muxOutConnector[34] = fifoOut[43][8];
              muxOutConnector[35] = fifoOut[44][8];
              muxOutConnector[36] = fifoOut[45][8];
              muxOutConnector[37] = fifoOut[46][8];
              muxOutConnector[38] = fifoOut[47][8];
              muxOutConnector[39] = fifoOut[48][8];
              muxOutConnector[40] = fifoOut[49][8];
              muxOutConnector[41] = fifoOut[50][8];
              muxOutConnector[42] = fifoOut[51][8];
              muxOutConnector[43] = fifoOut[26][7];
              muxOutConnector[44] = fifoOut[27][7];
              muxOutConnector[45] = fifoOut[28][7];
              muxOutConnector[46] = fifoOut[29][7];
              muxOutConnector[47] = fifoOut[30][7];
              muxOutConnector[48] = fifoOut[31][7];
              muxOutConnector[49] = fifoOut[32][7];
              muxOutConnector[50] = fifoOut[33][7];
              muxOutConnector[51] = fifoOut[34][7];
       end
       2: begin
              muxOutConnector[0] = fifoOut[44][3];
              muxOutConnector[1] = fifoOut[45][3];
              muxOutConnector[2] = fifoOut[46][3];
              muxOutConnector[3] = fifoOut[47][3];
              muxOutConnector[4] = fifoOut[48][3];
              muxOutConnector[5] = fifoOut[49][3];
              muxOutConnector[6] = fifoOut[50][3];
              muxOutConnector[7] = fifoOut[51][3];
              muxOutConnector[8] = fifoOut[26][2];
              muxOutConnector[9] = fifoOut[27][2];
              muxOutConnector[10] = fifoOut[28][2];
              muxOutConnector[11] = fifoOut[29][2];
              muxOutConnector[12] = fifoOut[30][2];
              muxOutConnector[13] = fifoOut[31][2];
              muxOutConnector[14] = fifoOut[32][2];
              muxOutConnector[15] = fifoOut[33][2];
              muxOutConnector[16] = fifoOut[34][2];
              muxOutConnector[17] = fifoOut[35][2];
              muxOutConnector[18] = fifoOut[36][2];
              muxOutConnector[19] = fifoOut[37][2];
              muxOutConnector[20] = fifoOut[38][2];
              muxOutConnector[21] = fifoOut[39][2];
              muxOutConnector[22] = fifoOut[40][2];
              muxOutConnector[23] = fifoOut[41][2];
              muxOutConnector[24] = fifoOut[42][2];
              muxOutConnector[25] = fifoOut[20][1];
              muxOutConnector[26] = fifoOut[35][8];
              muxOutConnector[27] = fifoOut[36][8];
              muxOutConnector[28] = fifoOut[37][8];
              muxOutConnector[29] = fifoOut[38][8];
              muxOutConnector[30] = fifoOut[39][8];
              muxOutConnector[31] = fifoOut[40][8];
              muxOutConnector[32] = fifoOut[41][8];
              muxOutConnector[33] = fifoOut[42][8];
              muxOutConnector[34] = fifoOut[43][8];
              muxOutConnector[35] = fifoOut[44][8];
              muxOutConnector[36] = fifoOut[45][8];
              muxOutConnector[37] = fifoOut[46][8];
              muxOutConnector[38] = fifoOut[47][8];
              muxOutConnector[39] = fifoOut[48][8];
              muxOutConnector[40] = fifoOut[49][8];
              muxOutConnector[41] = fifoOut[50][8];
              muxOutConnector[42] = fifoOut[51][8];
              muxOutConnector[43] = fifoOut[26][7];
              muxOutConnector[44] = fifoOut[27][7];
              muxOutConnector[45] = fifoOut[28][7];
              muxOutConnector[46] = fifoOut[29][7];
              muxOutConnector[47] = fifoOut[30][7];
              muxOutConnector[48] = fifoOut[31][7];
              muxOutConnector[49] = fifoOut[32][7];
              muxOutConnector[50] = fifoOut[33][7];
              muxOutConnector[51] = fifoOut[34][7];
       end
       3: begin
              muxOutConnector[0] = fifoOut[21][2];
              muxOutConnector[1] = fifoOut[22][2];
              muxOutConnector[2] = fifoOut[23][2];
              muxOutConnector[3] = fifoOut[24][2];
              muxOutConnector[4] = fifoOut[25][2];
              muxOutConnector[5] = fifoOut[0][1];
              muxOutConnector[6] = fifoOut[1][1];
              muxOutConnector[7] = fifoOut[2][1];
              muxOutConnector[8] = fifoOut[3][1];
              muxOutConnector[9] = fifoOut[4][1];
              muxOutConnector[10] = fifoOut[5][1];
              muxOutConnector[11] = fifoOut[6][1];
              muxOutConnector[12] = fifoOut[7][1];
              muxOutConnector[13] = fifoOut[8][1];
              muxOutConnector[14] = fifoOut[9][1];
              muxOutConnector[15] = fifoOut[10][1];
              muxOutConnector[16] = fifoOut[11][1];
              muxOutConnector[17] = fifoOut[12][1];
              muxOutConnector[18] = fifoOut[13][1];
              muxOutConnector[19] = fifoOut[14][1];
              muxOutConnector[20] = fifoOut[15][1];
              muxOutConnector[21] = fifoOut[16][1];
              muxOutConnector[22] = fifoOut[17][1];
              muxOutConnector[23] = fifoOut[18][1];
              muxOutConnector[24] = fifoOut[19][1];
              muxOutConnector[25] = fifoOut[20][1];
              muxOutConnector[26] = fifoOut[35][8];
              muxOutConnector[27] = fifoOut[36][8];
              muxOutConnector[28] = fifoOut[37][8];
              muxOutConnector[29] = fifoOut[38][8];
              muxOutConnector[30] = fifoOut[39][8];
              muxOutConnector[31] = fifoOut[40][8];
              muxOutConnector[32] = fifoOut[41][8];
              muxOutConnector[33] = fifoOut[42][8];
              muxOutConnector[34] = fifoOut[43][8];
              muxOutConnector[35] = fifoOut[44][8];
              muxOutConnector[36] = fifoOut[45][8];
              muxOutConnector[37] = fifoOut[46][8];
              muxOutConnector[38] = fifoOut[47][8];
              muxOutConnector[39] = fifoOut[48][8];
              muxOutConnector[40] = fifoOut[49][8];
              muxOutConnector[41] = fifoOut[50][8];
              muxOutConnector[42] = fifoOut[51][8];
              muxOutConnector[43] = fifoOut[26][7];
              muxOutConnector[44] = fifoOut[27][7];
              muxOutConnector[45] = fifoOut[28][7];
              muxOutConnector[46] = fifoOut[29][7];
              muxOutConnector[47] = fifoOut[30][7];
              muxOutConnector[48] = fifoOut[31][7];
              muxOutConnector[49] = fifoOut[32][7];
              muxOutConnector[50] = fifoOut[33][7];
              muxOutConnector[51] = fifoOut[34][7];
       end
       4: begin
              muxOutConnector[0] = fifoOut[21][2];
              muxOutConnector[1] = fifoOut[22][2];
              muxOutConnector[2] = fifoOut[23][2];
              muxOutConnector[3] = fifoOut[24][2];
              muxOutConnector[4] = fifoOut[25][2];
              muxOutConnector[5] = fifoOut[0][1];
              muxOutConnector[6] = fifoOut[1][1];
              muxOutConnector[7] = fifoOut[2][1];
              muxOutConnector[8] = fifoOut[3][1];
              muxOutConnector[9] = fifoOut[4][1];
              muxOutConnector[10] = fifoOut[5][1];
              muxOutConnector[11] = fifoOut[6][1];
              muxOutConnector[12] = fifoOut[7][1];
              muxOutConnector[13] = fifoOut[8][1];
              muxOutConnector[14] = fifoOut[9][1];
              muxOutConnector[15] = fifoOut[10][1];
              muxOutConnector[16] = fifoOut[11][1];
              muxOutConnector[17] = fifoOut[12][1];
              muxOutConnector[18] = fifoOut[13][1];
              muxOutConnector[19] = fifoOut[14][1];
              muxOutConnector[20] = fifoOut[15][1];
              muxOutConnector[21] = fifoOut[16][1];
              muxOutConnector[22] = fifoOut[17][1];
              muxOutConnector[23] = fifoOut[18][1];
              muxOutConnector[24] = fifoOut[19][1];
              muxOutConnector[25] = fifoOut[20][1];
              muxOutConnector[26] = fifoOut[35][8];
              muxOutConnector[27] = fifoOut[36][8];
              muxOutConnector[28] = fifoOut[37][8];
              muxOutConnector[29] = fifoOut[38][8];
              muxOutConnector[30] = fifoOut[39][8];
              muxOutConnector[31] = fifoOut[40][8];
              muxOutConnector[32] = fifoOut[41][8];
              muxOutConnector[33] = fifoOut[42][8];
              muxOutConnector[34] = fifoOut[43][8];
              muxOutConnector[35] = fifoOut[44][8];
              muxOutConnector[36] = fifoOut[45][8];
              muxOutConnector[37] = fifoOut[46][8];
              muxOutConnector[38] = fifoOut[47][8];
              muxOutConnector[39] = fifoOut[48][8];
              muxOutConnector[40] = fifoOut[49][8];
              muxOutConnector[41] = fifoOut[50][8];
              muxOutConnector[42] = fifoOut[51][8];
              muxOutConnector[43] = fifoOut[26][7];
              muxOutConnector[44] = fifoOut[27][7];
              muxOutConnector[45] = fifoOut[28][7];
              muxOutConnector[46] = fifoOut[29][7];
              muxOutConnector[47] = fifoOut[30][7];
              muxOutConnector[48] = fifoOut[31][7];
              muxOutConnector[49] = fifoOut[32][7];
              muxOutConnector[50] = fifoOut[33][7];
              muxOutConnector[51] = fifoOut[34][7];
       end
       5: begin
              muxOutConnector[0] = fifoOut[21][2];
              muxOutConnector[1] = fifoOut[22][2];
              muxOutConnector[2] = fifoOut[23][2];
              muxOutConnector[3] = fifoOut[24][2];
              muxOutConnector[4] = fifoOut[25][2];
              muxOutConnector[5] = fifoOut[0][1];
              muxOutConnector[6] = fifoOut[1][1];
              muxOutConnector[7] = fifoOut[2][1];
              muxOutConnector[8] = fifoOut[3][1];
              muxOutConnector[9] = fifoOut[4][1];
              muxOutConnector[10] = fifoOut[5][1];
              muxOutConnector[11] = fifoOut[6][1];
              muxOutConnector[12] = fifoOut[7][1];
              muxOutConnector[13] = fifoOut[8][1];
              muxOutConnector[14] = fifoOut[9][1];
              muxOutConnector[15] = fifoOut[10][1];
              muxOutConnector[16] = fifoOut[11][1];
              muxOutConnector[17] = fifoOut[12][1];
              muxOutConnector[18] = fifoOut[13][1];
              muxOutConnector[19] = fifoOut[14][1];
              muxOutConnector[20] = fifoOut[15][1];
              muxOutConnector[21] = fifoOut[16][1];
              muxOutConnector[22] = fifoOut[17][1];
              muxOutConnector[23] = fifoOut[18][1];
              muxOutConnector[24] = fifoOut[19][1];
              muxOutConnector[25] = fifoOut[20][1];
              muxOutConnector[26] = fifoOut[35][8];
              muxOutConnector[27] = fifoOut[36][8];
              muxOutConnector[28] = fifoOut[37][8];
              muxOutConnector[29] = fifoOut[38][8];
              muxOutConnector[30] = fifoOut[39][8];
              muxOutConnector[31] = fifoOut[40][8];
              muxOutConnector[32] = fifoOut[41][8];
              muxOutConnector[33] = fifoOut[42][8];
              muxOutConnector[34] = fifoOut[43][8];
              muxOutConnector[35] = fifoOut[44][8];
              muxOutConnector[36] = fifoOut[45][8];
              muxOutConnector[37] = fifoOut[46][8];
              muxOutConnector[38] = fifoOut[47][8];
              muxOutConnector[39] = fifoOut[48][8];
              muxOutConnector[40] = fifoOut[49][8];
              muxOutConnector[41] = fifoOut[50][8];
              muxOutConnector[42] = fifoOut[51][8];
              muxOutConnector[43] = fifoOut[26][7];
              muxOutConnector[44] = fifoOut[27][7];
              muxOutConnector[45] = fifoOut[28][7];
              muxOutConnector[46] = fifoOut[29][7];
              muxOutConnector[47] = fifoOut[30][7];
              muxOutConnector[48] = fifoOut[31][7];
              muxOutConnector[49] = fifoOut[32][7];
              muxOutConnector[50] = fifoOut[33][7];
              muxOutConnector[51] = fifoOut[34][7];
       end
       6: begin
              muxOutConnector[0] = fifoOut[21][2];
              muxOutConnector[1] = fifoOut[22][2];
              muxOutConnector[2] = fifoOut[23][2];
              muxOutConnector[3] = fifoOut[24][2];
              muxOutConnector[4] = fifoOut[25][2];
              muxOutConnector[5] = fifoOut[0][1];
              muxOutConnector[6] = fifoOut[1][1];
              muxOutConnector[7] = fifoOut[2][1];
              muxOutConnector[8] = fifoOut[3][1];
              muxOutConnector[9] = fifoOut[4][1];
              muxOutConnector[10] = fifoOut[5][1];
              muxOutConnector[11] = fifoOut[6][1];
              muxOutConnector[12] = fifoOut[7][1];
              muxOutConnector[13] = fifoOut[8][1];
              muxOutConnector[14] = fifoOut[9][1];
              muxOutConnector[15] = fifoOut[10][1];
              muxOutConnector[16] = fifoOut[11][1];
              muxOutConnector[17] = fifoOut[12][1];
              muxOutConnector[18] = fifoOut[13][1];
              muxOutConnector[19] = fifoOut[14][1];
              muxOutConnector[20] = fifoOut[15][1];
              muxOutConnector[21] = fifoOut[16][1];
              muxOutConnector[22] = fifoOut[17][1];
              muxOutConnector[23] = fifoOut[18][1];
              muxOutConnector[24] = fifoOut[19][1];
              muxOutConnector[25] = fifoOut[20][1];
              muxOutConnector[26] = fifoOut[35][8];
              muxOutConnector[27] = fifoOut[36][8];
              muxOutConnector[28] = fifoOut[37][8];
              muxOutConnector[29] = fifoOut[38][8];
              muxOutConnector[30] = fifoOut[39][8];
              muxOutConnector[31] = fifoOut[40][8];
              muxOutConnector[32] = fifoOut[41][8];
              muxOutConnector[33] = fifoOut[42][8];
              muxOutConnector[34] = fifoOut[43][8];
              muxOutConnector[35] = fifoOut[44][8];
              muxOutConnector[36] = fifoOut[45][8];
              muxOutConnector[37] = fifoOut[46][8];
              muxOutConnector[38] = fifoOut[47][8];
              muxOutConnector[39] = fifoOut[48][8];
              muxOutConnector[40] = fifoOut[49][8];
              muxOutConnector[41] = fifoOut[50][8];
              muxOutConnector[42] = fifoOut[51][8];
              muxOutConnector[43] = fifoOut[26][7];
              muxOutConnector[44] = fifoOut[27][7];
              muxOutConnector[45] = fifoOut[28][7];
              muxOutConnector[46] = fifoOut[29][7];
              muxOutConnector[47] = fifoOut[30][7];
              muxOutConnector[48] = fifoOut[31][7];
              muxOutConnector[49] = fifoOut[32][7];
              muxOutConnector[50] = fifoOut[33][7];
              muxOutConnector[51] = fifoOut[34][7];
       end
       7: begin
              muxOutConnector[0] = fifoOut[21][2];
              muxOutConnector[1] = fifoOut[22][2];
              muxOutConnector[2] = fifoOut[23][2];
              muxOutConnector[3] = fifoOut[24][2];
              muxOutConnector[4] = fifoOut[25][2];
              muxOutConnector[5] = fifoOut[0][1];
              muxOutConnector[6] = fifoOut[1][1];
              muxOutConnector[7] = fifoOut[2][1];
              muxOutConnector[8] = fifoOut[3][1];
              muxOutConnector[9] = fifoOut[4][1];
              muxOutConnector[10] = fifoOut[5][1];
              muxOutConnector[11] = fifoOut[6][1];
              muxOutConnector[12] = fifoOut[7][1];
              muxOutConnector[13] = fifoOut[8][1];
              muxOutConnector[14] = fifoOut[9][1];
              muxOutConnector[15] = fifoOut[10][1];
              muxOutConnector[16] = fifoOut[11][1];
              muxOutConnector[17] = fifoOut[12][1];
              muxOutConnector[18] = fifoOut[13][1];
              muxOutConnector[19] = fifoOut[14][1];
              muxOutConnector[20] = fifoOut[15][1];
              muxOutConnector[21] = fifoOut[16][1];
              muxOutConnector[22] = fifoOut[17][1];
              muxOutConnector[23] = fifoOut[18][1];
              muxOutConnector[24] = fifoOut[19][1];
              muxOutConnector[25] = fifoOut[20][1];
              muxOutConnector[26] = fifoOut[35][8];
              muxOutConnector[27] = fifoOut[36][8];
              muxOutConnector[28] = fifoOut[37][8];
              muxOutConnector[29] = fifoOut[38][8];
              muxOutConnector[30] = fifoOut[39][8];
              muxOutConnector[31] = fifoOut[40][8];
              muxOutConnector[32] = fifoOut[41][8];
              muxOutConnector[33] = fifoOut[42][8];
              muxOutConnector[34] = fifoOut[43][8];
              muxOutConnector[35] = fifoOut[44][8];
              muxOutConnector[36] = fifoOut[45][8];
              muxOutConnector[37] = fifoOut[46][8];
              muxOutConnector[38] = fifoOut[47][8];
              muxOutConnector[39] = fifoOut[48][8];
              muxOutConnector[40] = fifoOut[49][8];
              muxOutConnector[41] = fifoOut[50][8];
              muxOutConnector[42] = fifoOut[51][8];
              muxOutConnector[43] = fifoOut[26][7];
              muxOutConnector[44] = fifoOut[27][7];
              muxOutConnector[45] = fifoOut[28][7];
              muxOutConnector[46] = fifoOut[29][7];
              muxOutConnector[47] = fifoOut[30][7];
              muxOutConnector[48] = fifoOut[31][7];
              muxOutConnector[49] = fifoOut[32][7];
              muxOutConnector[50] = fifoOut[33][7];
              muxOutConnector[51] = fifoOut[34][7];
       end
       8: begin
              muxOutConnector[0] = fifoOut[21][2];
              muxOutConnector[1] = fifoOut[22][2];
              muxOutConnector[2] = fifoOut[23][2];
              muxOutConnector[3] = fifoOut[24][2];
              muxOutConnector[4] = fifoOut[25][2];
              muxOutConnector[5] = fifoOut[0][1];
              muxOutConnector[6] = fifoOut[1][1];
              muxOutConnector[7] = fifoOut[2][1];
              muxOutConnector[8] = fifoOut[3][1];
              muxOutConnector[9] = fifoOut[4][1];
              muxOutConnector[10] = fifoOut[5][1];
              muxOutConnector[11] = fifoOut[6][1];
              muxOutConnector[12] = fifoOut[7][1];
              muxOutConnector[13] = fifoOut[8][1];
              muxOutConnector[14] = fifoOut[9][1];
              muxOutConnector[15] = fifoOut[10][1];
              muxOutConnector[16] = fifoOut[11][1];
              muxOutConnector[17] = fifoOut[12][1];
              muxOutConnector[18] = fifoOut[13][1];
              muxOutConnector[19] = fifoOut[14][1];
              muxOutConnector[20] = fifoOut[15][1];
              muxOutConnector[21] = fifoOut[16][1];
              muxOutConnector[22] = fifoOut[17][1];
              muxOutConnector[23] = fifoOut[18][1];
              muxOutConnector[24] = fifoOut[19][1];
              muxOutConnector[25] = fifoOut[26][7];
              muxOutConnector[26] = fifoOut[35][8];
              muxOutConnector[27] = fifoOut[36][8];
              muxOutConnector[28] = fifoOut[37][8];
              muxOutConnector[29] = fifoOut[38][8];
              muxOutConnector[30] = fifoOut[39][8];
              muxOutConnector[31] = fifoOut[40][8];
              muxOutConnector[32] = fifoOut[41][8];
              muxOutConnector[33] = fifoOut[42][8];
              muxOutConnector[34] = fifoOut[20][7];
              muxOutConnector[35] = fifoOut[21][7];
              muxOutConnector[36] = fifoOut[22][7];
              muxOutConnector[37] = fifoOut[23][7];
              muxOutConnector[38] = fifoOut[24][7];
              muxOutConnector[39] = fifoOut[25][7];
              muxOutConnector[40] = fifoOut[0][6];
              muxOutConnector[41] = fifoOut[1][6];
              muxOutConnector[42] = fifoOut[2][6];
              muxOutConnector[43] = fifoOut[3][6];
              muxOutConnector[44] = fifoOut[4][6];
              muxOutConnector[45] = fifoOut[5][6];
              muxOutConnector[46] = fifoOut[6][6];
              muxOutConnector[47] = fifoOut[7][6];
              muxOutConnector[48] = fifoOut[8][6];
              muxOutConnector[49] = fifoOut[9][6];
              muxOutConnector[50] = fifoOut[10][6];
              muxOutConnector[51] = fifoOut[11][6];
       end
       9: begin
              muxOutConnector[0] = fifoOut[27][8];
              muxOutConnector[1] = fifoOut[28][8];
              muxOutConnector[2] = fifoOut[29][8];
              muxOutConnector[3] = fifoOut[30][8];
              muxOutConnector[4] = fifoOut[31][8];
              muxOutConnector[5] = fifoOut[32][8];
              muxOutConnector[6] = fifoOut[33][8];
              muxOutConnector[7] = fifoOut[34][8];
              muxOutConnector[8] = fifoOut[35][8];
              muxOutConnector[9] = fifoOut[36][8];
              muxOutConnector[10] = fifoOut[37][8];
              muxOutConnector[11] = fifoOut[38][8];
              muxOutConnector[12] = fifoOut[39][8];
              muxOutConnector[13] = fifoOut[40][8];
              muxOutConnector[14] = fifoOut[41][8];
              muxOutConnector[15] = fifoOut[42][8];
              muxOutConnector[16] = fifoOut[43][8];
              muxOutConnector[17] = fifoOut[44][8];
              muxOutConnector[18] = fifoOut[45][8];
              muxOutConnector[19] = fifoOut[46][8];
              muxOutConnector[20] = fifoOut[47][8];
              muxOutConnector[21] = fifoOut[48][8];
              muxOutConnector[22] = fifoOut[49][8];
              muxOutConnector[23] = fifoOut[50][8];
              muxOutConnector[24] = fifoOut[51][8];
              muxOutConnector[25] = fifoOut[26][7];
              muxOutConnector[26] = fifoOut[12][7];
              muxOutConnector[27] = fifoOut[13][7];
              muxOutConnector[28] = fifoOut[14][7];
              muxOutConnector[29] = fifoOut[15][7];
              muxOutConnector[30] = fifoOut[16][7];
              muxOutConnector[31] = fifoOut[17][7];
              muxOutConnector[32] = fifoOut[18][7];
              muxOutConnector[33] = fifoOut[19][7];
              muxOutConnector[34] = fifoOut[20][7];
              muxOutConnector[35] = fifoOut[21][7];
              muxOutConnector[36] = fifoOut[22][7];
              muxOutConnector[37] = fifoOut[23][7];
              muxOutConnector[38] = fifoOut[24][7];
              muxOutConnector[39] = fifoOut[25][7];
              muxOutConnector[40] = fifoOut[0][6];
              muxOutConnector[41] = fifoOut[1][6];
              muxOutConnector[42] = fifoOut[2][6];
              muxOutConnector[43] = fifoOut[3][6];
              muxOutConnector[44] = fifoOut[4][6];
              muxOutConnector[45] = fifoOut[5][6];
              muxOutConnector[46] = fifoOut[6][6];
              muxOutConnector[47] = fifoOut[7][6];
              muxOutConnector[48] = fifoOut[8][6];
              muxOutConnector[49] = fifoOut[9][6];
              muxOutConnector[50] = fifoOut[10][6];
              muxOutConnector[51] = fifoOut[11][6];
       end
       10: begin
              muxOutConnector[0] = fifoOut[27][8];
              muxOutConnector[1] = fifoOut[28][8];
              muxOutConnector[2] = fifoOut[29][8];
              muxOutConnector[3] = fifoOut[30][8];
              muxOutConnector[4] = fifoOut[31][8];
              muxOutConnector[5] = fifoOut[32][8];
              muxOutConnector[6] = fifoOut[33][8];
              muxOutConnector[7] = fifoOut[34][8];
              muxOutConnector[8] = fifoOut[35][8];
              muxOutConnector[9] = fifoOut[36][8];
              muxOutConnector[10] = fifoOut[37][8];
              muxOutConnector[11] = fifoOut[38][8];
              muxOutConnector[12] = fifoOut[39][8];
              muxOutConnector[13] = fifoOut[40][8];
              muxOutConnector[14] = fifoOut[41][8];
              muxOutConnector[15] = fifoOut[42][8];
              muxOutConnector[16] = fifoOut[43][8];
              muxOutConnector[17] = fifoOut[44][8];
              muxOutConnector[18] = fifoOut[45][8];
              muxOutConnector[19] = fifoOut[46][8];
              muxOutConnector[20] = fifoOut[47][8];
              muxOutConnector[21] = fifoOut[48][8];
              muxOutConnector[22] = fifoOut[49][8];
              muxOutConnector[23] = fifoOut[50][8];
              muxOutConnector[24] = fifoOut[51][8];
              muxOutConnector[25] = fifoOut[26][7];
              muxOutConnector[26] = fifoOut[12][7];
              muxOutConnector[27] = fifoOut[13][7];
              muxOutConnector[28] = fifoOut[14][7];
              muxOutConnector[29] = fifoOut[15][7];
              muxOutConnector[30] = fifoOut[16][7];
              muxOutConnector[31] = fifoOut[17][7];
              muxOutConnector[32] = fifoOut[18][7];
              muxOutConnector[33] = fifoOut[19][7];
              muxOutConnector[34] = fifoOut[20][7];
              muxOutConnector[35] = fifoOut[21][7];
              muxOutConnector[36] = fifoOut[22][7];
              muxOutConnector[37] = fifoOut[23][7];
              muxOutConnector[38] = fifoOut[24][7];
              muxOutConnector[39] = fifoOut[25][7];
              muxOutConnector[40] = fifoOut[0][6];
              muxOutConnector[41] = fifoOut[1][6];
              muxOutConnector[42] = fifoOut[2][6];
              muxOutConnector[43] = fifoOut[3][6];
              muxOutConnector[44] = fifoOut[4][6];
              muxOutConnector[45] = fifoOut[5][6];
              muxOutConnector[46] = fifoOut[6][6];
              muxOutConnector[47] = fifoOut[7][6];
              muxOutConnector[48] = fifoOut[8][6];
              muxOutConnector[49] = fifoOut[9][6];
              muxOutConnector[50] = fifoOut[10][6];
              muxOutConnector[51] = fifoOut[11][6];
       end
       11: begin
              muxOutConnector[0] = fifoOut[27][8];
              muxOutConnector[1] = fifoOut[28][8];
              muxOutConnector[2] = fifoOut[29][8];
              muxOutConnector[3] = fifoOut[30][8];
              muxOutConnector[4] = fifoOut[31][8];
              muxOutConnector[5] = fifoOut[32][8];
              muxOutConnector[6] = fifoOut[33][8];
              muxOutConnector[7] = fifoOut[34][8];
              muxOutConnector[8] = fifoOut[35][8];
              muxOutConnector[9] = fifoOut[36][8];
              muxOutConnector[10] = fifoOut[37][8];
              muxOutConnector[11] = fifoOut[38][8];
              muxOutConnector[12] = fifoOut[39][8];
              muxOutConnector[13] = fifoOut[40][8];
              muxOutConnector[14] = fifoOut[41][8];
              muxOutConnector[15] = fifoOut[42][8];
              muxOutConnector[16] = fifoOut[43][8];
              muxOutConnector[17] = fifoOut[44][8];
              muxOutConnector[18] = fifoOut[45][8];
              muxOutConnector[19] = fifoOut[46][8];
              muxOutConnector[20] = fifoOut[47][8];
              muxOutConnector[21] = fifoOut[48][8];
              muxOutConnector[22] = fifoOut[49][8];
              muxOutConnector[23] = fifoOut[50][8];
              muxOutConnector[24] = fifoOut[51][8];
              muxOutConnector[25] = fifoOut[26][7];
              muxOutConnector[26] = fifoOut[12][7];
              muxOutConnector[27] = fifoOut[13][7];
              muxOutConnector[28] = fifoOut[14][7];
              muxOutConnector[29] = fifoOut[15][7];
              muxOutConnector[30] = fifoOut[16][7];
              muxOutConnector[31] = fifoOut[17][7];
              muxOutConnector[32] = fifoOut[18][7];
              muxOutConnector[33] = fifoOut[19][7];
              muxOutConnector[34] = fifoOut[20][7];
              muxOutConnector[35] = fifoOut[21][7];
              muxOutConnector[36] = fifoOut[22][7];
              muxOutConnector[37] = fifoOut[23][7];
              muxOutConnector[38] = fifoOut[24][7];
              muxOutConnector[39] = fifoOut[25][7];
              muxOutConnector[40] = fifoOut[0][6];
              muxOutConnector[41] = fifoOut[1][6];
              muxOutConnector[42] = fifoOut[2][6];
              muxOutConnector[43] = fifoOut[3][6];
              muxOutConnector[44] = fifoOut[4][6];
              muxOutConnector[45] = fifoOut[5][6];
              muxOutConnector[46] = fifoOut[6][6];
              muxOutConnector[47] = fifoOut[7][6];
              muxOutConnector[48] = fifoOut[8][6];
              muxOutConnector[49] = fifoOut[9][6];
              muxOutConnector[50] = fifoOut[10][6];
              muxOutConnector[51] = fifoOut[11][6];
       end
       12: begin
              muxOutConnector[0] = fifoOut[27][8];
              muxOutConnector[1] = fifoOut[28][8];
              muxOutConnector[2] = fifoOut[29][8];
              muxOutConnector[3] = fifoOut[30][8];
              muxOutConnector[4] = fifoOut[31][8];
              muxOutConnector[5] = fifoOut[32][8];
              muxOutConnector[6] = fifoOut[33][8];
              muxOutConnector[7] = fifoOut[34][8];
              muxOutConnector[8] = fifoOut[35][8];
              muxOutConnector[9] = fifoOut[36][8];
              muxOutConnector[10] = fifoOut[37][8];
              muxOutConnector[11] = fifoOut[38][8];
              muxOutConnector[12] = fifoOut[39][8];
              muxOutConnector[13] = fifoOut[40][8];
              muxOutConnector[14] = fifoOut[41][8];
              muxOutConnector[15] = fifoOut[42][8];
              muxOutConnector[16] = fifoOut[43][8];
              muxOutConnector[17] = fifoOut[44][8];
              muxOutConnector[18] = fifoOut[45][8];
              muxOutConnector[19] = fifoOut[46][8];
              muxOutConnector[20] = fifoOut[47][8];
              muxOutConnector[21] = fifoOut[48][8];
              muxOutConnector[22] = fifoOut[49][8];
              muxOutConnector[23] = fifoOut[50][8];
              muxOutConnector[24] = fifoOut[51][8];
              muxOutConnector[25] = fifoOut[26][7];
              muxOutConnector[26] = fifoOut[12][7];
              muxOutConnector[27] = fifoOut[13][7];
              muxOutConnector[28] = fifoOut[14][7];
              muxOutConnector[29] = fifoOut[15][7];
              muxOutConnector[30] = fifoOut[16][7];
              muxOutConnector[31] = fifoOut[17][7];
              muxOutConnector[32] = fifoOut[18][7];
              muxOutConnector[33] = fifoOut[19][7];
              muxOutConnector[34] = fifoOut[20][7];
              muxOutConnector[35] = fifoOut[21][7];
              muxOutConnector[36] = fifoOut[22][7];
              muxOutConnector[37] = fifoOut[23][7];
              muxOutConnector[38] = fifoOut[24][7];
              muxOutConnector[39] = fifoOut[25][7];
              muxOutConnector[40] = fifoOut[0][6];
              muxOutConnector[41] = fifoOut[1][6];
              muxOutConnector[42] = fifoOut[2][6];
              muxOutConnector[43] = fifoOut[3][6];
              muxOutConnector[44] = fifoOut[4][6];
              muxOutConnector[45] = fifoOut[5][6];
              muxOutConnector[46] = fifoOut[6][6];
              muxOutConnector[47] = fifoOut[7][6];
              muxOutConnector[48] = fifoOut[8][6];
              muxOutConnector[49] = fifoOut[9][6];
              muxOutConnector[50] = fifoOut[10][6];
              muxOutConnector[51] = fifoOut[11][6];
       end
       13: begin
              muxOutConnector[0] = fifoOut[27][8];
              muxOutConnector[1] = fifoOut[28][8];
              muxOutConnector[2] = fifoOut[29][8];
              muxOutConnector[3] = fifoOut[30][8];
              muxOutConnector[4] = fifoOut[31][8];
              muxOutConnector[5] = fifoOut[32][8];
              muxOutConnector[6] = fifoOut[33][8];
              muxOutConnector[7] = fifoOut[34][8];
              muxOutConnector[8] = fifoOut[35][8];
              muxOutConnector[9] = fifoOut[36][8];
              muxOutConnector[10] = fifoOut[37][8];
              muxOutConnector[11] = fifoOut[38][8];
              muxOutConnector[12] = fifoOut[39][8];
              muxOutConnector[13] = fifoOut[40][8];
              muxOutConnector[14] = fifoOut[41][8];
              muxOutConnector[15] = fifoOut[42][8];
              muxOutConnector[16] = fifoOut[43][8];
              muxOutConnector[17] = fifoOut[44][8];
              muxOutConnector[18] = fifoOut[45][8];
              muxOutConnector[19] = fifoOut[46][8];
              muxOutConnector[20] = fifoOut[47][8];
              muxOutConnector[21] = fifoOut[48][8];
              muxOutConnector[22] = fifoOut[49][8];
              muxOutConnector[23] = fifoOut[50][8];
              muxOutConnector[24] = fifoOut[51][8];
              muxOutConnector[25] = fifoOut[26][7];
              muxOutConnector[26] = fifoOut[12][7];
              muxOutConnector[27] = fifoOut[13][7];
              muxOutConnector[28] = fifoOut[14][7];
              muxOutConnector[29] = fifoOut[15][7];
              muxOutConnector[30] = fifoOut[16][7];
              muxOutConnector[31] = fifoOut[17][7];
              muxOutConnector[32] = fifoOut[18][7];
              muxOutConnector[33] = fifoOut[19][7];
              muxOutConnector[34] = fifoOut[20][7];
              muxOutConnector[35] = fifoOut[21][7];
              muxOutConnector[36] = fifoOut[22][7];
              muxOutConnector[37] = fifoOut[23][7];
              muxOutConnector[38] = fifoOut[24][7];
              muxOutConnector[39] = fifoOut[25][7];
              muxOutConnector[40] = fifoOut[0][6];
              muxOutConnector[41] = fifoOut[1][6];
              muxOutConnector[42] = fifoOut[2][6];
              muxOutConnector[43] = fifoOut[3][6];
              muxOutConnector[44] = fifoOut[4][6];
              muxOutConnector[45] = fifoOut[5][6];
              muxOutConnector[46] = fifoOut[6][6];
              muxOutConnector[47] = fifoOut[7][6];
              muxOutConnector[48] = fifoOut[8][6];
              muxOutConnector[49] = fifoOut[9][6];
              muxOutConnector[50] = fifoOut[10][6];
              muxOutConnector[51] = fifoOut[11][6];
       end
       14: begin
              muxOutConnector[0] = fifoOut[27][8];
              muxOutConnector[1] = fifoOut[28][8];
              muxOutConnector[2] = fifoOut[29][8];
              muxOutConnector[3] = fifoOut[30][8];
              muxOutConnector[4] = fifoOut[31][8];
              muxOutConnector[5] = fifoOut[32][8];
              muxOutConnector[6] = fifoOut[33][8];
              muxOutConnector[7] = fifoOut[34][8];
              muxOutConnector[8] = fifoOut[35][8];
              muxOutConnector[9] = fifoOut[36][8];
              muxOutConnector[10] = fifoOut[37][8];
              muxOutConnector[11] = fifoOut[38][8];
              muxOutConnector[12] = fifoOut[39][8];
              muxOutConnector[13] = fifoOut[40][8];
              muxOutConnector[14] = fifoOut[41][8];
              muxOutConnector[15] = fifoOut[42][8];
              muxOutConnector[16] = fifoOut[43][8];
              muxOutConnector[17] = fifoOut[44][8];
              muxOutConnector[18] = fifoOut[45][8];
              muxOutConnector[19] = fifoOut[46][8];
              muxOutConnector[20] = fifoOut[47][8];
              muxOutConnector[21] = fifoOut[48][8];
              muxOutConnector[22] = fifoOut[49][8];
              muxOutConnector[23] = fifoOut[50][8];
              muxOutConnector[24] = fifoOut[51][8];
              muxOutConnector[25] = fifoOut[26][7];
              muxOutConnector[26] = fifoOut[12][7];
              muxOutConnector[27] = fifoOut[13][7];
              muxOutConnector[28] = fifoOut[14][7];
              muxOutConnector[29] = fifoOut[15][7];
              muxOutConnector[30] = fifoOut[16][7];
              muxOutConnector[31] = fifoOut[17][7];
              muxOutConnector[32] = fifoOut[18][7];
              muxOutConnector[33] = fifoOut[19][7];
              muxOutConnector[34] = fifoOut[26][13];
              muxOutConnector[35] = fifoOut[27][13];
              muxOutConnector[36] = fifoOut[28][13];
              muxOutConnector[37] = fifoOut[29][13];
              muxOutConnector[38] = fifoOut[30][13];
              muxOutConnector[39] = fifoOut[31][13];
              muxOutConnector[40] = fifoOut[32][13];
              muxOutConnector[41] = fifoOut[33][13];
              muxOutConnector[42] = fifoOut[34][13];
              muxOutConnector[43] = fifoOut[35][13];
              muxOutConnector[44] = fifoOut[36][13];
              muxOutConnector[45] = fifoOut[37][13];
              muxOutConnector[46] = fifoOut[38][13];
              muxOutConnector[47] = fifoOut[39][13];
              muxOutConnector[48] = fifoOut[40][13];
              muxOutConnector[49] = fifoOut[41][13];
              muxOutConnector[50] = fifoOut[42][13];
              muxOutConnector[51] = fifoOut[43][13];
       end
       15: begin
              muxOutConnector[0] = fifoOut[27][8];
              muxOutConnector[1] = fifoOut[28][8];
              muxOutConnector[2] = fifoOut[29][8];
              muxOutConnector[3] = fifoOut[30][8];
              muxOutConnector[4] = fifoOut[31][8];
              muxOutConnector[5] = fifoOut[32][8];
              muxOutConnector[6] = fifoOut[33][8];
              muxOutConnector[7] = fifoOut[34][8];
              muxOutConnector[8] = fifoOut[35][8];
              muxOutConnector[9] = fifoOut[36][8];
              muxOutConnector[10] = fifoOut[37][8];
              muxOutConnector[11] = fifoOut[38][8];
              muxOutConnector[12] = fifoOut[39][8];
              muxOutConnector[13] = fifoOut[40][8];
              muxOutConnector[14] = fifoOut[41][8];
              muxOutConnector[15] = fifoOut[42][8];
              muxOutConnector[16] = fifoOut[43][8];
              muxOutConnector[17] = fifoOut[44][8];
              muxOutConnector[18] = fifoOut[45][8];
              muxOutConnector[19] = fifoOut[46][8];
              muxOutConnector[20] = fifoOut[47][8];
              muxOutConnector[21] = fifoOut[48][8];
              muxOutConnector[22] = fifoOut[49][8];
              muxOutConnector[23] = fifoOut[50][8];
              muxOutConnector[24] = fifoOut[51][8];
              muxOutConnector[25] = fifoOut[26][7];
              muxOutConnector[26] = fifoOut[12][7];
              muxOutConnector[27] = fifoOut[13][7];
              muxOutConnector[28] = fifoOut[14][7];
              muxOutConnector[29] = fifoOut[15][7];
              muxOutConnector[30] = fifoOut[16][7];
              muxOutConnector[31] = fifoOut[17][7];
              muxOutConnector[32] = fifoOut[18][7];
              muxOutConnector[33] = fifoOut[19][7];
              muxOutConnector[34] = fifoOut[26][13];
              muxOutConnector[35] = fifoOut[27][13];
              muxOutConnector[36] = fifoOut[28][13];
              muxOutConnector[37] = fifoOut[29][13];
              muxOutConnector[38] = fifoOut[30][13];
              muxOutConnector[39] = fifoOut[31][13];
              muxOutConnector[40] = fifoOut[32][13];
              muxOutConnector[41] = fifoOut[33][13];
              muxOutConnector[42] = fifoOut[34][13];
              muxOutConnector[43] = fifoOut[35][13];
              muxOutConnector[44] = fifoOut[36][13];
              muxOutConnector[45] = fifoOut[37][13];
              muxOutConnector[46] = fifoOut[38][13];
              muxOutConnector[47] = fifoOut[39][13];
              muxOutConnector[48] = fifoOut[40][13];
              muxOutConnector[49] = fifoOut[41][13];
              muxOutConnector[50] = fifoOut[42][13];
              muxOutConnector[51] = fifoOut[43][13];
       end
       16: begin
              muxOutConnector[0] = fifoOut[27][8];
              muxOutConnector[1] = fifoOut[28][8];
              muxOutConnector[2] = fifoOut[29][8];
              muxOutConnector[3] = fifoOut[30][8];
              muxOutConnector[4] = fifoOut[31][8];
              muxOutConnector[5] = fifoOut[32][8];
              muxOutConnector[6] = fifoOut[33][8];
              muxOutConnector[7] = fifoOut[34][8];
              muxOutConnector[8] = fifoOut[35][8];
              muxOutConnector[9] = fifoOut[36][8];
              muxOutConnector[10] = fifoOut[37][8];
              muxOutConnector[11] = fifoOut[38][8];
              muxOutConnector[12] = fifoOut[39][8];
              muxOutConnector[13] = fifoOut[40][8];
              muxOutConnector[14] = fifoOut[41][8];
              muxOutConnector[15] = fifoOut[42][8];
              muxOutConnector[16] = fifoOut[43][8];
              muxOutConnector[17] = fifoOut[44][8];
              muxOutConnector[18] = fifoOut[45][8];
              muxOutConnector[19] = fifoOut[46][8];
              muxOutConnector[20] = fifoOut[47][8];
              muxOutConnector[21] = fifoOut[48][8];
              muxOutConnector[22] = fifoOut[49][8];
              muxOutConnector[23] = fifoOut[50][8];
              muxOutConnector[24] = fifoOut[51][8];
              muxOutConnector[25] = fifoOut[26][7];
              muxOutConnector[26] = fifoOut[12][7];
              muxOutConnector[27] = fifoOut[13][7];
              muxOutConnector[28] = fifoOut[14][7];
              muxOutConnector[29] = fifoOut[15][7];
              muxOutConnector[30] = fifoOut[16][7];
              muxOutConnector[31] = fifoOut[17][7];
              muxOutConnector[32] = fifoOut[18][7];
              muxOutConnector[33] = fifoOut[19][7];
              muxOutConnector[34] = fifoOut[26][13];
              muxOutConnector[35] = fifoOut[27][13];
              muxOutConnector[36] = fifoOut[28][13];
              muxOutConnector[37] = fifoOut[29][13];
              muxOutConnector[38] = fifoOut[30][13];
              muxOutConnector[39] = fifoOut[31][13];
              muxOutConnector[40] = fifoOut[32][13];
              muxOutConnector[41] = fifoOut[33][13];
              muxOutConnector[42] = fifoOut[34][13];
              muxOutConnector[43] = fifoOut[35][13];
              muxOutConnector[44] = fifoOut[36][13];
              muxOutConnector[45] = fifoOut[37][13];
              muxOutConnector[46] = fifoOut[38][13];
              muxOutConnector[47] = fifoOut[39][13];
              muxOutConnector[48] = fifoOut[40][13];
              muxOutConnector[49] = fifoOut[41][13];
              muxOutConnector[50] = fifoOut[42][13];
              muxOutConnector[51] = fifoOut[43][13];
       end
       17: begin
              muxOutConnector[0] = fifoOut[27][8];
              muxOutConnector[1] = fifoOut[28][8];
              muxOutConnector[2] = fifoOut[29][8];
              muxOutConnector[3] = fifoOut[30][8];
              muxOutConnector[4] = fifoOut[31][8];
              muxOutConnector[5] = fifoOut[32][8];
              muxOutConnector[6] = fifoOut[33][8];
              muxOutConnector[7] = fifoOut[34][8];
              muxOutConnector[8] = fifoOut[35][8];
              muxOutConnector[9] = fifoOut[36][8];
              muxOutConnector[10] = fifoOut[37][8];
              muxOutConnector[11] = fifoOut[38][8];
              muxOutConnector[12] = fifoOut[39][8];
              muxOutConnector[13] = fifoOut[40][8];
              muxOutConnector[14] = fifoOut[41][8];
              muxOutConnector[15] = fifoOut[42][8];
              muxOutConnector[16] = fifoOut[43][8];
              muxOutConnector[17] = fifoOut[44][8];
              muxOutConnector[18] = fifoOut[45][8];
              muxOutConnector[19] = fifoOut[46][8];
              muxOutConnector[20] = fifoOut[47][8];
              muxOutConnector[21] = fifoOut[48][8];
              muxOutConnector[22] = fifoOut[49][8];
              muxOutConnector[23] = fifoOut[50][8];
              muxOutConnector[24] = fifoOut[51][8];
              muxOutConnector[25] = fifoOut[26][7];
              muxOutConnector[26] = fifoOut[12][7];
              muxOutConnector[27] = fifoOut[13][7];
              muxOutConnector[28] = fifoOut[14][7];
              muxOutConnector[29] = fifoOut[15][7];
              muxOutConnector[30] = fifoOut[16][7];
              muxOutConnector[31] = fifoOut[17][7];
              muxOutConnector[32] = fifoOut[18][7];
              muxOutConnector[33] = fifoOut[19][7];
              muxOutConnector[34] = fifoOut[26][13];
              muxOutConnector[35] = fifoOut[27][13];
              muxOutConnector[36] = fifoOut[28][13];
              muxOutConnector[37] = fifoOut[29][13];
              muxOutConnector[38] = fifoOut[30][13];
              muxOutConnector[39] = fifoOut[31][13];
              muxOutConnector[40] = fifoOut[32][13];
              muxOutConnector[41] = fifoOut[33][13];
              muxOutConnector[42] = fifoOut[34][13];
              muxOutConnector[43] = fifoOut[35][13];
              muxOutConnector[44] = fifoOut[36][13];
              muxOutConnector[45] = fifoOut[37][13];
              muxOutConnector[46] = fifoOut[38][13];
              muxOutConnector[47] = fifoOut[39][13];
              muxOutConnector[48] = fifoOut[40][13];
              muxOutConnector[49] = fifoOut[41][13];
              muxOutConnector[50] = fifoOut[42][13];
              muxOutConnector[51] = fifoOut[43][13];
       end
       18: begin
              muxOutConnector[0] = fifoOut[27][8];
              muxOutConnector[1] = fifoOut[28][8];
              muxOutConnector[2] = fifoOut[29][8];
              muxOutConnector[3] = fifoOut[30][8];
              muxOutConnector[4] = fifoOut[31][8];
              muxOutConnector[5] = fifoOut[32][8];
              muxOutConnector[6] = fifoOut[33][8];
              muxOutConnector[7] = fifoOut[34][8];
              muxOutConnector[8] = fifoOut[35][8];
              muxOutConnector[9] = fifoOut[36][8];
              muxOutConnector[10] = fifoOut[37][8];
              muxOutConnector[11] = fifoOut[38][8];
              muxOutConnector[12] = fifoOut[39][8];
              muxOutConnector[13] = fifoOut[40][8];
              muxOutConnector[14] = fifoOut[41][8];
              muxOutConnector[15] = fifoOut[42][8];
              muxOutConnector[16] = fifoOut[43][8];
              muxOutConnector[17] = fifoOut[44][8];
              muxOutConnector[18] = fifoOut[45][8];
              muxOutConnector[19] = fifoOut[46][8];
              muxOutConnector[20] = fifoOut[47][8];
              muxOutConnector[21] = fifoOut[48][8];
              muxOutConnector[22] = fifoOut[49][8];
              muxOutConnector[23] = fifoOut[50][8];
              muxOutConnector[24] = fifoOut[51][8];
              muxOutConnector[25] = fifoOut[26][7];
              muxOutConnector[26] = fifoOut[12][7];
              muxOutConnector[27] = fifoOut[13][7];
              muxOutConnector[28] = fifoOut[14][7];
              muxOutConnector[29] = fifoOut[15][7];
              muxOutConnector[30] = fifoOut[16][7];
              muxOutConnector[31] = fifoOut[17][7];
              muxOutConnector[32] = fifoOut[18][7];
              muxOutConnector[33] = fifoOut[19][7];
              muxOutConnector[34] = fifoOut[26][13];
              muxOutConnector[35] = fifoOut[27][13];
              muxOutConnector[36] = fifoOut[28][13];
              muxOutConnector[37] = fifoOut[29][13];
              muxOutConnector[38] = fifoOut[30][13];
              muxOutConnector[39] = fifoOut[31][13];
              muxOutConnector[40] = fifoOut[32][13];
              muxOutConnector[41] = fifoOut[33][13];
              muxOutConnector[42] = fifoOut[34][13];
              muxOutConnector[43] = fifoOut[35][13];
              muxOutConnector[44] = fifoOut[36][13];
              muxOutConnector[45] = fifoOut[37][13];
              muxOutConnector[46] = fifoOut[38][13];
              muxOutConnector[47] = fifoOut[39][13];
              muxOutConnector[48] = fifoOut[40][13];
              muxOutConnector[49] = fifoOut[41][13];
              muxOutConnector[50] = fifoOut[42][13];
              muxOutConnector[51] = fifoOut[43][13];
       end
       19: begin
              muxOutConnector[0] = fifoOut[27][8];
              muxOutConnector[1] = fifoOut[28][8];
              muxOutConnector[2] = fifoOut[29][8];
              muxOutConnector[3] = fifoOut[30][8];
              muxOutConnector[4] = fifoOut[31][8];
              muxOutConnector[5] = fifoOut[32][8];
              muxOutConnector[6] = fifoOut[33][8];
              muxOutConnector[7] = fifoOut[34][8];
              muxOutConnector[8] = fifoOut[35][8];
              muxOutConnector[9] = fifoOut[36][8];
              muxOutConnector[10] = fifoOut[37][8];
              muxOutConnector[11] = fifoOut[38][8];
              muxOutConnector[12] = fifoOut[39][8];
              muxOutConnector[13] = fifoOut[40][8];
              muxOutConnector[14] = fifoOut[41][8];
              muxOutConnector[15] = fifoOut[42][8];
              muxOutConnector[16] = fifoOut[43][8];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[12][7];
              muxOutConnector[27] = fifoOut[13][7];
              muxOutConnector[28] = fifoOut[14][7];
              muxOutConnector[29] = fifoOut[15][7];
              muxOutConnector[30] = fifoOut[16][7];
              muxOutConnector[31] = fifoOut[17][7];
              muxOutConnector[32] = fifoOut[18][7];
              muxOutConnector[33] = fifoOut[19][7];
              muxOutConnector[34] = fifoOut[26][13];
              muxOutConnector[35] = fifoOut[27][13];
              muxOutConnector[36] = fifoOut[28][13];
              muxOutConnector[37] = fifoOut[29][13];
              muxOutConnector[38] = fifoOut[30][13];
              muxOutConnector[39] = fifoOut[31][13];
              muxOutConnector[40] = fifoOut[32][13];
              muxOutConnector[41] = fifoOut[33][13];
              muxOutConnector[42] = fifoOut[34][13];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
