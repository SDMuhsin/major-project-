`timescale 1ns / 1ps
module LMem0To1_511_circ5_ys_scripted(
        muxOut,
        ly0In,
        wr_en,
        feedback_en,
        rd_address,
        rd_en,
        clk,
        rst
);
input feedback_en;
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 11;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        if(feedback_en) begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= fifoOut[i][c-1];
         end
        end
        else begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= ly0InConnector[i];
         end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[46][5];
              muxOutConnector[1] = fifoOut[47][5];
              muxOutConnector[2] = fifoOut[48][5];
              muxOutConnector[3] = fifoOut[49][5];
              muxOutConnector[4] = fifoOut[50][5];
              muxOutConnector[5] = fifoOut[51][5];
              muxOutConnector[6] = fifoOut[26][4];
              muxOutConnector[7] = fifoOut[27][4];
              muxOutConnector[8] = fifoOut[28][4];
              muxOutConnector[9] = fifoOut[29][4];
              muxOutConnector[10] = fifoOut[30][4];
              muxOutConnector[11] = fifoOut[31][4];
              muxOutConnector[12] = fifoOut[32][4];
              muxOutConnector[13] = fifoOut[33][4];
              muxOutConnector[14] = fifoOut[34][4];
              muxOutConnector[15] = fifoOut[35][4];
              muxOutConnector[16] = fifoOut[36][4];
              muxOutConnector[17] = fifoOut[37][4];
              muxOutConnector[18] = fifoOut[38][4];
              muxOutConnector[19] = fifoOut[39][4];
              muxOutConnector[20] = fifoOut[40][4];
              muxOutConnector[21] = fifoOut[41][4];
              muxOutConnector[22] = fifoOut[42][4];
              muxOutConnector[23] = fifoOut[43][4];
              muxOutConnector[24] = fifoOut[44][4];
              muxOutConnector[25] = fifoOut[45][4];
              muxOutConnector[26] = fifoOut[18][7];
              muxOutConnector[27] = fifoOut[19][7];
              muxOutConnector[28] = fifoOut[20][7];
              muxOutConnector[29] = fifoOut[21][7];
              muxOutConnector[30] = fifoOut[22][7];
              muxOutConnector[31] = fifoOut[23][7];
              muxOutConnector[32] = fifoOut[24][7];
              muxOutConnector[33] = fifoOut[25][7];
              muxOutConnector[34] = fifoOut[0][6];
              muxOutConnector[35] = fifoOut[1][6];
              muxOutConnector[36] = fifoOut[2][6];
              muxOutConnector[37] = fifoOut[3][6];
              muxOutConnector[38] = fifoOut[4][6];
              muxOutConnector[39] = fifoOut[5][6];
              muxOutConnector[40] = fifoOut[6][6];
              muxOutConnector[41] = fifoOut[7][6];
              muxOutConnector[42] = fifoOut[8][6];
              muxOutConnector[43] = fifoOut[9][6];
              muxOutConnector[44] = fifoOut[10][6];
              muxOutConnector[45] = fifoOut[11][6];
              muxOutConnector[46] = fifoOut[12][6];
              muxOutConnector[47] = fifoOut[13][6];
              muxOutConnector[48] = fifoOut[14][6];
              muxOutConnector[49] = fifoOut[15][6];
              muxOutConnector[50] = fifoOut[16][6];
              muxOutConnector[51] = fifoOut[17][6];
       end
       1: begin
              muxOutConnector[0] = fifoOut[46][5];
              muxOutConnector[1] = fifoOut[47][5];
              muxOutConnector[2] = fifoOut[48][5];
              muxOutConnector[3] = fifoOut[49][5];
              muxOutConnector[4] = fifoOut[50][5];
              muxOutConnector[5] = fifoOut[51][5];
              muxOutConnector[6] = fifoOut[26][4];
              muxOutConnector[7] = fifoOut[27][4];
              muxOutConnector[8] = fifoOut[28][4];
              muxOutConnector[9] = fifoOut[29][4];
              muxOutConnector[10] = fifoOut[30][4];
              muxOutConnector[11] = fifoOut[31][4];
              muxOutConnector[12] = fifoOut[32][4];
              muxOutConnector[13] = fifoOut[33][4];
              muxOutConnector[14] = fifoOut[34][4];
              muxOutConnector[15] = fifoOut[35][4];
              muxOutConnector[16] = fifoOut[36][4];
              muxOutConnector[17] = fifoOut[37][4];
              muxOutConnector[18] = fifoOut[38][4];
              muxOutConnector[19] = fifoOut[39][4];
              muxOutConnector[20] = fifoOut[40][4];
              muxOutConnector[21] = fifoOut[41][4];
              muxOutConnector[22] = fifoOut[42][4];
              muxOutConnector[23] = fifoOut[43][4];
              muxOutConnector[24] = fifoOut[44][4];
              muxOutConnector[25] = fifoOut[45][4];
              muxOutConnector[26] = fifoOut[18][7];
              muxOutConnector[27] = fifoOut[19][7];
              muxOutConnector[28] = fifoOut[20][7];
              muxOutConnector[29] = fifoOut[21][7];
              muxOutConnector[30] = fifoOut[22][7];
              muxOutConnector[31] = fifoOut[23][7];
              muxOutConnector[32] = fifoOut[24][7];
              muxOutConnector[33] = fifoOut[25][7];
              muxOutConnector[34] = fifoOut[0][6];
              muxOutConnector[35] = fifoOut[1][6];
              muxOutConnector[36] = fifoOut[2][6];
              muxOutConnector[37] = fifoOut[3][6];
              muxOutConnector[38] = fifoOut[4][6];
              muxOutConnector[39] = fifoOut[5][6];
              muxOutConnector[40] = fifoOut[6][6];
              muxOutConnector[41] = fifoOut[7][6];
              muxOutConnector[42] = fifoOut[8][6];
              muxOutConnector[43] = fifoOut[9][6];
              muxOutConnector[44] = fifoOut[10][6];
              muxOutConnector[45] = fifoOut[11][6];
              muxOutConnector[46] = fifoOut[12][6];
              muxOutConnector[47] = fifoOut[13][6];
              muxOutConnector[48] = fifoOut[14][6];
              muxOutConnector[49] = fifoOut[15][6];
              muxOutConnector[50] = fifoOut[16][6];
              muxOutConnector[51] = fifoOut[17][6];
       end
       2: begin
              muxOutConnector[0] = fifoOut[46][5];
              muxOutConnector[1] = fifoOut[47][5];
              muxOutConnector[2] = fifoOut[48][5];
              muxOutConnector[3] = fifoOut[49][5];
              muxOutConnector[4] = fifoOut[50][5];
              muxOutConnector[5] = fifoOut[51][5];
              muxOutConnector[6] = fifoOut[26][4];
              muxOutConnector[7] = fifoOut[27][4];
              muxOutConnector[8] = fifoOut[28][4];
              muxOutConnector[9] = fifoOut[29][4];
              muxOutConnector[10] = fifoOut[30][4];
              muxOutConnector[11] = fifoOut[31][4];
              muxOutConnector[12] = fifoOut[32][4];
              muxOutConnector[13] = fifoOut[33][4];
              muxOutConnector[14] = fifoOut[34][4];
              muxOutConnector[15] = fifoOut[35][4];
              muxOutConnector[16] = fifoOut[36][4];
              muxOutConnector[17] = fifoOut[37][4];
              muxOutConnector[18] = fifoOut[38][4];
              muxOutConnector[19] = fifoOut[39][4];
              muxOutConnector[20] = fifoOut[40][4];
              muxOutConnector[21] = fifoOut[41][4];
              muxOutConnector[22] = fifoOut[42][4];
              muxOutConnector[23] = fifoOut[43][4];
              muxOutConnector[24] = fifoOut[44][4];
              muxOutConnector[25] = fifoOut[45][4];
              muxOutConnector[26] = fifoOut[18][7];
              muxOutConnector[27] = fifoOut[19][7];
              muxOutConnector[28] = fifoOut[20][7];
              muxOutConnector[29] = fifoOut[21][7];
              muxOutConnector[30] = fifoOut[22][7];
              muxOutConnector[31] = fifoOut[23][7];
              muxOutConnector[32] = fifoOut[24][7];
              muxOutConnector[33] = fifoOut[25][7];
              muxOutConnector[34] = fifoOut[0][6];
              muxOutConnector[35] = fifoOut[1][6];
              muxOutConnector[36] = fifoOut[2][6];
              muxOutConnector[37] = fifoOut[3][6];
              muxOutConnector[38] = fifoOut[4][6];
              muxOutConnector[39] = fifoOut[5][6];
              muxOutConnector[40] = fifoOut[6][6];
              muxOutConnector[41] = fifoOut[7][6];
              muxOutConnector[42] = fifoOut[8][6];
              muxOutConnector[43] = fifoOut[9][6];
              muxOutConnector[44] = fifoOut[10][6];
              muxOutConnector[45] = fifoOut[11][6];
              muxOutConnector[46] = fifoOut[12][6];
              muxOutConnector[47] = fifoOut[13][6];
              muxOutConnector[48] = fifoOut[14][6];
              muxOutConnector[49] = fifoOut[15][6];
              muxOutConnector[50] = fifoOut[16][6];
              muxOutConnector[51] = fifoOut[17][6];
       end
       3: begin
              muxOutConnector[0] = fifoOut[46][5];
              muxOutConnector[1] = fifoOut[47][5];
              muxOutConnector[2] = fifoOut[48][5];
              muxOutConnector[3] = fifoOut[49][5];
              muxOutConnector[4] = fifoOut[50][5];
              muxOutConnector[5] = fifoOut[51][5];
              muxOutConnector[6] = fifoOut[26][4];
              muxOutConnector[7] = fifoOut[27][4];
              muxOutConnector[8] = fifoOut[28][4];
              muxOutConnector[9] = fifoOut[29][4];
              muxOutConnector[10] = fifoOut[30][4];
              muxOutConnector[11] = fifoOut[31][4];
              muxOutConnector[12] = fifoOut[32][4];
              muxOutConnector[13] = fifoOut[33][4];
              muxOutConnector[14] = fifoOut[34][4];
              muxOutConnector[15] = fifoOut[35][4];
              muxOutConnector[16] = fifoOut[36][4];
              muxOutConnector[17] = fifoOut[37][4];
              muxOutConnector[18] = fifoOut[38][4];
              muxOutConnector[19] = fifoOut[39][4];
              muxOutConnector[20] = fifoOut[40][4];
              muxOutConnector[21] = fifoOut[41][4];
              muxOutConnector[22] = fifoOut[42][4];
              muxOutConnector[23] = fifoOut[43][4];
              muxOutConnector[24] = fifoOut[44][4];
              muxOutConnector[25] = fifoOut[45][4];
              muxOutConnector[26] = fifoOut[18][7];
              muxOutConnector[27] = fifoOut[19][7];
              muxOutConnector[28] = fifoOut[20][7];
              muxOutConnector[29] = fifoOut[21][7];
              muxOutConnector[30] = fifoOut[22][7];
              muxOutConnector[31] = fifoOut[23][7];
              muxOutConnector[32] = fifoOut[24][7];
              muxOutConnector[33] = fifoOut[25][7];
              muxOutConnector[34] = fifoOut[0][6];
              muxOutConnector[35] = fifoOut[1][6];
              muxOutConnector[36] = fifoOut[2][6];
              muxOutConnector[37] = fifoOut[3][6];
              muxOutConnector[38] = fifoOut[4][6];
              muxOutConnector[39] = fifoOut[5][6];
              muxOutConnector[40] = fifoOut[6][6];
              muxOutConnector[41] = fifoOut[7][6];
              muxOutConnector[42] = fifoOut[8][6];
              muxOutConnector[43] = fifoOut[9][6];
              muxOutConnector[44] = fifoOut[10][6];
              muxOutConnector[45] = fifoOut[11][6];
              muxOutConnector[46] = fifoOut[12][6];
              muxOutConnector[47] = fifoOut[13][6];
              muxOutConnector[48] = fifoOut[14][6];
              muxOutConnector[49] = fifoOut[15][6];
              muxOutConnector[50] = fifoOut[16][6];
              muxOutConnector[51] = fifoOut[17][6];
       end
       4: begin
              muxOutConnector[0] = fifoOut[46][5];
              muxOutConnector[1] = fifoOut[47][5];
              muxOutConnector[2] = fifoOut[48][5];
              muxOutConnector[3] = fifoOut[49][5];
              muxOutConnector[4] = fifoOut[50][5];
              muxOutConnector[5] = fifoOut[51][5];
              muxOutConnector[6] = fifoOut[26][4];
              muxOutConnector[7] = fifoOut[27][4];
              muxOutConnector[8] = fifoOut[28][4];
              muxOutConnector[9] = fifoOut[29][4];
              muxOutConnector[10] = fifoOut[30][4];
              muxOutConnector[11] = fifoOut[31][4];
              muxOutConnector[12] = fifoOut[32][4];
              muxOutConnector[13] = fifoOut[33][4];
              muxOutConnector[14] = fifoOut[34][4];
              muxOutConnector[15] = fifoOut[35][4];
              muxOutConnector[16] = fifoOut[36][4];
              muxOutConnector[17] = fifoOut[37][4];
              muxOutConnector[18] = fifoOut[38][4];
              muxOutConnector[19] = fifoOut[39][4];
              muxOutConnector[20] = fifoOut[40][4];
              muxOutConnector[21] = fifoOut[41][4];
              muxOutConnector[22] = fifoOut[42][4];
              muxOutConnector[23] = fifoOut[24][3];
              muxOutConnector[24] = fifoOut[25][3];
              muxOutConnector[25] = fifoOut[0][2];
              muxOutConnector[26] = fifoOut[18][7];
              muxOutConnector[27] = fifoOut[19][7];
              muxOutConnector[28] = fifoOut[20][7];
              muxOutConnector[29] = fifoOut[21][7];
              muxOutConnector[30] = fifoOut[22][7];
              muxOutConnector[31] = fifoOut[23][7];
              muxOutConnector[32] = fifoOut[24][7];
              muxOutConnector[33] = fifoOut[25][7];
              muxOutConnector[34] = fifoOut[0][6];
              muxOutConnector[35] = fifoOut[1][6];
              muxOutConnector[36] = fifoOut[2][6];
              muxOutConnector[37] = fifoOut[3][6];
              muxOutConnector[38] = fifoOut[4][6];
              muxOutConnector[39] = fifoOut[5][6];
              muxOutConnector[40] = fifoOut[6][6];
              muxOutConnector[41] = fifoOut[7][6];
              muxOutConnector[42] = fifoOut[8][6];
              muxOutConnector[43] = fifoOut[9][6];
              muxOutConnector[44] = fifoOut[10][6];
              muxOutConnector[45] = fifoOut[11][6];
              muxOutConnector[46] = fifoOut[12][6];
              muxOutConnector[47] = fifoOut[13][6];
              muxOutConnector[48] = fifoOut[14][6];
              muxOutConnector[49] = fifoOut[15][6];
              muxOutConnector[50] = fifoOut[16][6];
              muxOutConnector[51] = fifoOut[17][6];
       end
       5: begin
              muxOutConnector[0] = fifoOut[1][3];
              muxOutConnector[1] = fifoOut[2][3];
              muxOutConnector[2] = fifoOut[3][3];
              muxOutConnector[3] = fifoOut[4][3];
              muxOutConnector[4] = fifoOut[5][3];
              muxOutConnector[5] = fifoOut[6][3];
              muxOutConnector[6] = fifoOut[7][3];
              muxOutConnector[7] = fifoOut[8][3];
              muxOutConnector[8] = fifoOut[9][3];
              muxOutConnector[9] = fifoOut[10][3];
              muxOutConnector[10] = fifoOut[11][3];
              muxOutConnector[11] = fifoOut[12][3];
              muxOutConnector[12] = fifoOut[13][3];
              muxOutConnector[13] = fifoOut[14][3];
              muxOutConnector[14] = fifoOut[15][3];
              muxOutConnector[15] = fifoOut[16][3];
              muxOutConnector[16] = fifoOut[17][3];
              muxOutConnector[17] = fifoOut[18][3];
              muxOutConnector[18] = fifoOut[19][3];
              muxOutConnector[19] = fifoOut[20][3];
              muxOutConnector[20] = fifoOut[21][3];
              muxOutConnector[21] = fifoOut[22][3];
              muxOutConnector[22] = fifoOut[23][3];
              muxOutConnector[23] = fifoOut[24][3];
              muxOutConnector[24] = fifoOut[25][3];
              muxOutConnector[25] = fifoOut[0][2];
              muxOutConnector[26] = fifoOut[18][7];
              muxOutConnector[27] = fifoOut[19][7];
              muxOutConnector[28] = fifoOut[20][7];
              muxOutConnector[29] = fifoOut[21][7];
              muxOutConnector[30] = fifoOut[22][7];
              muxOutConnector[31] = fifoOut[23][7];
              muxOutConnector[32] = fifoOut[24][7];
              muxOutConnector[33] = fifoOut[25][7];
              muxOutConnector[34] = fifoOut[0][6];
              muxOutConnector[35] = fifoOut[1][6];
              muxOutConnector[36] = fifoOut[2][6];
              muxOutConnector[37] = fifoOut[3][6];
              muxOutConnector[38] = fifoOut[4][6];
              muxOutConnector[39] = fifoOut[5][6];
              muxOutConnector[40] = fifoOut[6][6];
              muxOutConnector[41] = fifoOut[7][6];
              muxOutConnector[42] = fifoOut[8][6];
              muxOutConnector[43] = fifoOut[9][6];
              muxOutConnector[44] = fifoOut[10][6];
              muxOutConnector[45] = fifoOut[11][6];
              muxOutConnector[46] = fifoOut[12][6];
              muxOutConnector[47] = fifoOut[13][6];
              muxOutConnector[48] = fifoOut[14][6];
              muxOutConnector[49] = fifoOut[15][6];
              muxOutConnector[50] = fifoOut[16][6];
              muxOutConnector[51] = fifoOut[17][6];
       end
       6: begin
              muxOutConnector[0] = fifoOut[1][3];
              muxOutConnector[1] = fifoOut[2][3];
              muxOutConnector[2] = fifoOut[3][3];
              muxOutConnector[3] = fifoOut[4][3];
              muxOutConnector[4] = fifoOut[5][3];
              muxOutConnector[5] = fifoOut[6][3];
              muxOutConnector[6] = fifoOut[7][3];
              muxOutConnector[7] = fifoOut[8][3];
              muxOutConnector[8] = fifoOut[9][3];
              muxOutConnector[9] = fifoOut[10][3];
              muxOutConnector[10] = fifoOut[11][3];
              muxOutConnector[11] = fifoOut[12][3];
              muxOutConnector[12] = fifoOut[13][3];
              muxOutConnector[13] = fifoOut[14][3];
              muxOutConnector[14] = fifoOut[15][3];
              muxOutConnector[15] = fifoOut[16][3];
              muxOutConnector[16] = fifoOut[17][3];
              muxOutConnector[17] = fifoOut[18][3];
              muxOutConnector[18] = fifoOut[19][3];
              muxOutConnector[19] = fifoOut[20][3];
              muxOutConnector[20] = fifoOut[21][3];
              muxOutConnector[21] = fifoOut[22][3];
              muxOutConnector[22] = fifoOut[23][3];
              muxOutConnector[23] = fifoOut[24][3];
              muxOutConnector[24] = fifoOut[25][3];
              muxOutConnector[25] = fifoOut[0][2];
              muxOutConnector[26] = fifoOut[18][7];
              muxOutConnector[27] = fifoOut[19][7];
              muxOutConnector[28] = fifoOut[20][7];
              muxOutConnector[29] = fifoOut[21][7];
              muxOutConnector[30] = fifoOut[22][7];
              muxOutConnector[31] = fifoOut[23][7];
              muxOutConnector[32] = fifoOut[24][7];
              muxOutConnector[33] = fifoOut[25][7];
              muxOutConnector[34] = fifoOut[0][6];
              muxOutConnector[35] = fifoOut[1][6];
              muxOutConnector[36] = fifoOut[2][6];
              muxOutConnector[37] = fifoOut[3][6];
              muxOutConnector[38] = fifoOut[4][6];
              muxOutConnector[39] = fifoOut[5][6];
              muxOutConnector[40] = fifoOut[6][6];
              muxOutConnector[41] = fifoOut[7][6];
              muxOutConnector[42] = fifoOut[8][6];
              muxOutConnector[43] = fifoOut[9][6];
              muxOutConnector[44] = fifoOut[10][6];
              muxOutConnector[45] = fifoOut[11][6];
              muxOutConnector[46] = fifoOut[12][6];
              muxOutConnector[47] = fifoOut[13][6];
              muxOutConnector[48] = fifoOut[14][6];
              muxOutConnector[49] = fifoOut[15][6];
              muxOutConnector[50] = fifoOut[16][6];
              muxOutConnector[51] = fifoOut[45][5];
       end
       7: begin
              muxOutConnector[0] = fifoOut[1][3];
              muxOutConnector[1] = fifoOut[2][3];
              muxOutConnector[2] = fifoOut[3][3];
              muxOutConnector[3] = fifoOut[4][3];
              muxOutConnector[4] = fifoOut[5][3];
              muxOutConnector[5] = fifoOut[6][3];
              muxOutConnector[6] = fifoOut[7][3];
              muxOutConnector[7] = fifoOut[8][3];
              muxOutConnector[8] = fifoOut[9][3];
              muxOutConnector[9] = fifoOut[10][3];
              muxOutConnector[10] = fifoOut[11][3];
              muxOutConnector[11] = fifoOut[12][3];
              muxOutConnector[12] = fifoOut[13][3];
              muxOutConnector[13] = fifoOut[14][3];
              muxOutConnector[14] = fifoOut[15][3];
              muxOutConnector[15] = fifoOut[16][3];
              muxOutConnector[16] = fifoOut[17][3];
              muxOutConnector[17] = fifoOut[18][3];
              muxOutConnector[18] = fifoOut[19][3];
              muxOutConnector[19] = fifoOut[20][3];
              muxOutConnector[20] = fifoOut[21][3];
              muxOutConnector[21] = fifoOut[22][3];
              muxOutConnector[22] = fifoOut[23][3];
              muxOutConnector[23] = fifoOut[24][3];
              muxOutConnector[24] = fifoOut[25][3];
              muxOutConnector[25] = fifoOut[0][2];
              muxOutConnector[26] = fifoOut[46][6];
              muxOutConnector[27] = fifoOut[47][6];
              muxOutConnector[28] = fifoOut[48][6];
              muxOutConnector[29] = fifoOut[49][6];
              muxOutConnector[30] = fifoOut[50][6];
              muxOutConnector[31] = fifoOut[51][6];
              muxOutConnector[32] = fifoOut[26][5];
              muxOutConnector[33] = fifoOut[27][5];
              muxOutConnector[34] = fifoOut[28][5];
              muxOutConnector[35] = fifoOut[29][5];
              muxOutConnector[36] = fifoOut[30][5];
              muxOutConnector[37] = fifoOut[31][5];
              muxOutConnector[38] = fifoOut[32][5];
              muxOutConnector[39] = fifoOut[33][5];
              muxOutConnector[40] = fifoOut[34][5];
              muxOutConnector[41] = fifoOut[35][5];
              muxOutConnector[42] = fifoOut[36][5];
              muxOutConnector[43] = fifoOut[37][5];
              muxOutConnector[44] = fifoOut[38][5];
              muxOutConnector[45] = fifoOut[39][5];
              muxOutConnector[46] = fifoOut[40][5];
              muxOutConnector[47] = fifoOut[41][5];
              muxOutConnector[48] = fifoOut[42][5];
              muxOutConnector[49] = fifoOut[43][5];
              muxOutConnector[50] = fifoOut[44][5];
              muxOutConnector[51] = fifoOut[45][5];
       end
       8: begin
              muxOutConnector[0] = fifoOut[1][3];
              muxOutConnector[1] = fifoOut[2][3];
              muxOutConnector[2] = fifoOut[3][3];
              muxOutConnector[3] = fifoOut[4][3];
              muxOutConnector[4] = fifoOut[5][3];
              muxOutConnector[5] = fifoOut[6][3];
              muxOutConnector[6] = fifoOut[7][3];
              muxOutConnector[7] = fifoOut[8][3];
              muxOutConnector[8] = fifoOut[9][3];
              muxOutConnector[9] = fifoOut[10][3];
              muxOutConnector[10] = fifoOut[11][3];
              muxOutConnector[11] = fifoOut[12][3];
              muxOutConnector[12] = fifoOut[13][3];
              muxOutConnector[13] = fifoOut[14][3];
              muxOutConnector[14] = fifoOut[15][3];
              muxOutConnector[15] = fifoOut[16][3];
              muxOutConnector[16] = fifoOut[17][3];
              muxOutConnector[17] = fifoOut[18][3];
              muxOutConnector[18] = fifoOut[19][3];
              muxOutConnector[19] = fifoOut[20][3];
              muxOutConnector[20] = fifoOut[21][3];
              muxOutConnector[21] = fifoOut[22][3];
              muxOutConnector[22] = fifoOut[23][3];
              muxOutConnector[23] = fifoOut[24][3];
              muxOutConnector[24] = fifoOut[25][3];
              muxOutConnector[25] = fifoOut[0][2];
              muxOutConnector[26] = fifoOut[46][6];
              muxOutConnector[27] = fifoOut[47][6];
              muxOutConnector[28] = fifoOut[48][6];
              muxOutConnector[29] = fifoOut[49][6];
              muxOutConnector[30] = fifoOut[50][6];
              muxOutConnector[31] = fifoOut[51][6];
              muxOutConnector[32] = fifoOut[26][5];
              muxOutConnector[33] = fifoOut[27][5];
              muxOutConnector[34] = fifoOut[28][5];
              muxOutConnector[35] = fifoOut[29][5];
              muxOutConnector[36] = fifoOut[30][5];
              muxOutConnector[37] = fifoOut[31][5];
              muxOutConnector[38] = fifoOut[32][5];
              muxOutConnector[39] = fifoOut[33][5];
              muxOutConnector[40] = fifoOut[34][5];
              muxOutConnector[41] = fifoOut[35][5];
              muxOutConnector[42] = fifoOut[36][5];
              muxOutConnector[43] = fifoOut[37][5];
              muxOutConnector[44] = fifoOut[38][5];
              muxOutConnector[45] = fifoOut[39][5];
              muxOutConnector[46] = fifoOut[40][5];
              muxOutConnector[47] = fifoOut[41][5];
              muxOutConnector[48] = fifoOut[42][5];
              muxOutConnector[49] = fifoOut[43][5];
              muxOutConnector[50] = fifoOut[44][5];
              muxOutConnector[51] = fifoOut[45][5];
       end
       9: begin
              muxOutConnector[0] = fifoOut[1][3];
              muxOutConnector[1] = fifoOut[2][3];
              muxOutConnector[2] = fifoOut[3][3];
              muxOutConnector[3] = fifoOut[4][3];
              muxOutConnector[4] = fifoOut[5][3];
              muxOutConnector[5] = fifoOut[6][3];
              muxOutConnector[6] = fifoOut[7][3];
              muxOutConnector[7] = fifoOut[8][3];
              muxOutConnector[8] = fifoOut[9][3];
              muxOutConnector[9] = fifoOut[10][3];
              muxOutConnector[10] = fifoOut[11][3];
              muxOutConnector[11] = fifoOut[12][3];
              muxOutConnector[12] = fifoOut[13][3];
              muxOutConnector[13] = fifoOut[14][3];
              muxOutConnector[14] = fifoOut[15][3];
              muxOutConnector[15] = fifoOut[16][3];
              muxOutConnector[16] = fifoOut[17][3];
              muxOutConnector[17] = fifoOut[18][3];
              muxOutConnector[18] = fifoOut[19][3];
              muxOutConnector[19] = fifoOut[20][3];
              muxOutConnector[20] = fifoOut[21][3];
              muxOutConnector[21] = fifoOut[22][3];
              muxOutConnector[22] = fifoOut[23][3];
              muxOutConnector[23] = fifoOut[24][3];
              muxOutConnector[24] = fifoOut[25][3];
              muxOutConnector[25] = fifoOut[0][2];
              muxOutConnector[26] = fifoOut[46][6];
              muxOutConnector[27] = fifoOut[47][6];
              muxOutConnector[28] = fifoOut[48][6];
              muxOutConnector[29] = fifoOut[49][6];
              muxOutConnector[30] = fifoOut[50][6];
              muxOutConnector[31] = fifoOut[51][6];
              muxOutConnector[32] = fifoOut[26][5];
              muxOutConnector[33] = fifoOut[27][5];
              muxOutConnector[34] = fifoOut[28][5];
              muxOutConnector[35] = fifoOut[29][5];
              muxOutConnector[36] = fifoOut[30][5];
              muxOutConnector[37] = fifoOut[31][5];
              muxOutConnector[38] = fifoOut[32][5];
              muxOutConnector[39] = fifoOut[33][5];
              muxOutConnector[40] = fifoOut[34][5];
              muxOutConnector[41] = fifoOut[35][5];
              muxOutConnector[42] = fifoOut[36][5];
              muxOutConnector[43] = fifoOut[37][5];
              muxOutConnector[44] = fifoOut[38][5];
              muxOutConnector[45] = fifoOut[39][5];
              muxOutConnector[46] = fifoOut[40][5];
              muxOutConnector[47] = fifoOut[41][5];
              muxOutConnector[48] = fifoOut[42][5];
              muxOutConnector[49] = fifoOut[43][5];
              muxOutConnector[50] = fifoOut[44][5];
              muxOutConnector[51] = fifoOut[45][5];
       end
       10: begin
              muxOutConnector[0] = fifoOut[1][3];
              muxOutConnector[1] = fifoOut[2][3];
              muxOutConnector[2] = fifoOut[3][3];
              muxOutConnector[3] = fifoOut[4][3];
              muxOutConnector[4] = fifoOut[5][3];
              muxOutConnector[5] = fifoOut[6][3];
              muxOutConnector[6] = fifoOut[7][3];
              muxOutConnector[7] = fifoOut[8][3];
              muxOutConnector[8] = fifoOut[9][3];
              muxOutConnector[9] = fifoOut[10][3];
              muxOutConnector[10] = fifoOut[11][3];
              muxOutConnector[11] = fifoOut[12][3];
              muxOutConnector[12] = fifoOut[13][3];
              muxOutConnector[13] = fifoOut[14][3];
              muxOutConnector[14] = fifoOut[15][3];
              muxOutConnector[15] = fifoOut[16][3];
              muxOutConnector[16] = fifoOut[17][3];
              muxOutConnector[17] = fifoOut[18][3];
              muxOutConnector[18] = fifoOut[19][3];
              muxOutConnector[19] = fifoOut[20][3];
              muxOutConnector[20] = fifoOut[21][3];
              muxOutConnector[21] = fifoOut[22][3];
              muxOutConnector[22] = fifoOut[23][3];
              muxOutConnector[23] = fifoOut[24][3];
              muxOutConnector[24] = fifoOut[25][3];
              muxOutConnector[25] = fifoOut[0][2];
              muxOutConnector[26] = fifoOut[46][6];
              muxOutConnector[27] = fifoOut[47][6];
              muxOutConnector[28] = fifoOut[48][6];
              muxOutConnector[29] = fifoOut[49][6];
              muxOutConnector[30] = fifoOut[50][6];
              muxOutConnector[31] = fifoOut[51][6];
              muxOutConnector[32] = fifoOut[26][5];
              muxOutConnector[33] = fifoOut[27][5];
              muxOutConnector[34] = fifoOut[28][5];
              muxOutConnector[35] = fifoOut[29][5];
              muxOutConnector[36] = fifoOut[30][5];
              muxOutConnector[37] = fifoOut[31][5];
              muxOutConnector[38] = fifoOut[32][5];
              muxOutConnector[39] = fifoOut[33][5];
              muxOutConnector[40] = fifoOut[34][5];
              muxOutConnector[41] = fifoOut[35][5];
              muxOutConnector[42] = fifoOut[36][5];
              muxOutConnector[43] = fifoOut[37][5];
              muxOutConnector[44] = fifoOut[38][5];
              muxOutConnector[45] = fifoOut[39][5];
              muxOutConnector[46] = fifoOut[40][5];
              muxOutConnector[47] = fifoOut[41][5];
              muxOutConnector[48] = fifoOut[42][5];
              muxOutConnector[49] = fifoOut[43][5];
              muxOutConnector[50] = fifoOut[44][5];
              muxOutConnector[51] = fifoOut[45][5];
       end
       11: begin
              muxOutConnector[0] = fifoOut[1][3];
              muxOutConnector[1] = fifoOut[2][3];
              muxOutConnector[2] = fifoOut[3][3];
              muxOutConnector[3] = fifoOut[4][3];
              muxOutConnector[4] = fifoOut[5][3];
              muxOutConnector[5] = fifoOut[6][3];
              muxOutConnector[6] = fifoOut[7][3];
              muxOutConnector[7] = fifoOut[8][3];
              muxOutConnector[8] = fifoOut[9][3];
              muxOutConnector[9] = fifoOut[10][3];
              muxOutConnector[10] = fifoOut[11][3];
              muxOutConnector[11] = fifoOut[12][3];
              muxOutConnector[12] = fifoOut[13][3];
              muxOutConnector[13] = fifoOut[14][3];
              muxOutConnector[14] = fifoOut[15][3];
              muxOutConnector[15] = fifoOut[16][3];
              muxOutConnector[16] = fifoOut[17][3];
              muxOutConnector[17] = fifoOut[18][3];
              muxOutConnector[18] = fifoOut[19][3];
              muxOutConnector[19] = fifoOut[20][3];
              muxOutConnector[20] = fifoOut[21][3];
              muxOutConnector[21] = fifoOut[22][3];
              muxOutConnector[22] = fifoOut[23][3];
              muxOutConnector[23] = fifoOut[24][3];
              muxOutConnector[24] = fifoOut[25][3];
              muxOutConnector[25] = fifoOut[0][2];
              muxOutConnector[26] = fifoOut[46][6];
              muxOutConnector[27] = fifoOut[47][6];
              muxOutConnector[28] = fifoOut[48][6];
              muxOutConnector[29] = fifoOut[49][6];
              muxOutConnector[30] = fifoOut[50][6];
              muxOutConnector[31] = fifoOut[51][6];
              muxOutConnector[32] = fifoOut[26][5];
              muxOutConnector[33] = fifoOut[27][5];
              muxOutConnector[34] = fifoOut[28][5];
              muxOutConnector[35] = fifoOut[29][5];
              muxOutConnector[36] = fifoOut[30][5];
              muxOutConnector[37] = fifoOut[31][5];
              muxOutConnector[38] = fifoOut[32][5];
              muxOutConnector[39] = fifoOut[33][5];
              muxOutConnector[40] = fifoOut[34][5];
              muxOutConnector[41] = fifoOut[35][5];
              muxOutConnector[42] = fifoOut[36][5];
              muxOutConnector[43] = fifoOut[37][5];
              muxOutConnector[44] = fifoOut[38][5];
              muxOutConnector[45] = fifoOut[39][5];
              muxOutConnector[46] = fifoOut[40][5];
              muxOutConnector[47] = fifoOut[41][5];
              muxOutConnector[48] = fifoOut[42][5];
              muxOutConnector[49] = fifoOut[43][5];
              muxOutConnector[50] = fifoOut[44][5];
              muxOutConnector[51] = fifoOut[45][5];
       end
       12: begin
              muxOutConnector[0] = fifoOut[1][3];
              muxOutConnector[1] = fifoOut[2][3];
              muxOutConnector[2] = fifoOut[3][3];
              muxOutConnector[3] = fifoOut[4][3];
              muxOutConnector[4] = fifoOut[5][3];
              muxOutConnector[5] = fifoOut[6][3];
              muxOutConnector[6] = fifoOut[7][3];
              muxOutConnector[7] = fifoOut[8][3];
              muxOutConnector[8] = fifoOut[9][3];
              muxOutConnector[9] = fifoOut[10][3];
              muxOutConnector[10] = fifoOut[11][3];
              muxOutConnector[11] = fifoOut[12][3];
              muxOutConnector[12] = fifoOut[13][3];
              muxOutConnector[13] = fifoOut[14][3];
              muxOutConnector[14] = fifoOut[15][3];
              muxOutConnector[15] = fifoOut[16][3];
              muxOutConnector[16] = fifoOut[17][3];
              muxOutConnector[17] = fifoOut[18][3];
              muxOutConnector[18] = fifoOut[19][3];
              muxOutConnector[19] = fifoOut[20][3];
              muxOutConnector[20] = fifoOut[21][3];
              muxOutConnector[21] = fifoOut[22][3];
              muxOutConnector[22] = fifoOut[23][3];
              muxOutConnector[23] = fifoOut[24][3];
              muxOutConnector[24] = fifoOut[25][3];
              muxOutConnector[25] = fifoOut[0][2];
              muxOutConnector[26] = fifoOut[46][6];
              muxOutConnector[27] = fifoOut[47][6];
              muxOutConnector[28] = fifoOut[48][6];
              muxOutConnector[29] = fifoOut[49][6];
              muxOutConnector[30] = fifoOut[50][6];
              muxOutConnector[31] = fifoOut[51][6];
              muxOutConnector[32] = fifoOut[26][5];
              muxOutConnector[33] = fifoOut[27][5];
              muxOutConnector[34] = fifoOut[28][5];
              muxOutConnector[35] = fifoOut[29][5];
              muxOutConnector[36] = fifoOut[30][5];
              muxOutConnector[37] = fifoOut[31][5];
              muxOutConnector[38] = fifoOut[32][5];
              muxOutConnector[39] = fifoOut[33][5];
              muxOutConnector[40] = fifoOut[34][5];
              muxOutConnector[41] = fifoOut[35][5];
              muxOutConnector[42] = fifoOut[36][5];
              muxOutConnector[43] = fifoOut[37][5];
              muxOutConnector[44] = fifoOut[38][5];
              muxOutConnector[45] = fifoOut[39][5];
              muxOutConnector[46] = fifoOut[40][5];
              muxOutConnector[47] = fifoOut[41][5];
              muxOutConnector[48] = fifoOut[42][5];
              muxOutConnector[49] = fifoOut[43][5];
              muxOutConnector[50] = fifoOut[44][5];
              muxOutConnector[51] = fifoOut[45][5];
       end
       13: begin
              muxOutConnector[0] = fifoOut[1][3];
              muxOutConnector[1] = fifoOut[2][3];
              muxOutConnector[2] = fifoOut[3][3];
              muxOutConnector[3] = fifoOut[4][3];
              muxOutConnector[4] = fifoOut[5][3];
              muxOutConnector[5] = fifoOut[6][3];
              muxOutConnector[6] = fifoOut[7][3];
              muxOutConnector[7] = fifoOut[8][3];
              muxOutConnector[8] = fifoOut[9][3];
              muxOutConnector[9] = fifoOut[10][3];
              muxOutConnector[10] = fifoOut[11][3];
              muxOutConnector[11] = fifoOut[12][3];
              muxOutConnector[12] = fifoOut[13][3];
              muxOutConnector[13] = fifoOut[14][3];
              muxOutConnector[14] = fifoOut[15][3];
              muxOutConnector[15] = fifoOut[16][3];
              muxOutConnector[16] = fifoOut[17][3];
              muxOutConnector[17] = fifoOut[18][3];
              muxOutConnector[18] = fifoOut[19][3];
              muxOutConnector[19] = fifoOut[20][3];
              muxOutConnector[20] = fifoOut[21][3];
              muxOutConnector[21] = fifoOut[22][3];
              muxOutConnector[22] = fifoOut[23][3];
              muxOutConnector[23] = fifoOut[24][3];
              muxOutConnector[24] = fifoOut[25][3];
              muxOutConnector[25] = fifoOut[0][2];
              muxOutConnector[26] = fifoOut[46][6];
              muxOutConnector[27] = fifoOut[47][6];
              muxOutConnector[28] = fifoOut[48][6];
              muxOutConnector[29] = fifoOut[49][6];
              muxOutConnector[30] = fifoOut[50][6];
              muxOutConnector[31] = fifoOut[51][6];
              muxOutConnector[32] = fifoOut[26][5];
              muxOutConnector[33] = fifoOut[27][5];
              muxOutConnector[34] = fifoOut[28][5];
              muxOutConnector[35] = fifoOut[29][5];
              muxOutConnector[36] = fifoOut[30][5];
              muxOutConnector[37] = fifoOut[31][5];
              muxOutConnector[38] = fifoOut[32][5];
              muxOutConnector[39] = fifoOut[33][5];
              muxOutConnector[40] = fifoOut[34][5];
              muxOutConnector[41] = fifoOut[35][5];
              muxOutConnector[42] = fifoOut[36][5];
              muxOutConnector[43] = fifoOut[37][5];
              muxOutConnector[44] = fifoOut[38][5];
              muxOutConnector[45] = fifoOut[39][5];
              muxOutConnector[46] = fifoOut[40][5];
              muxOutConnector[47] = fifoOut[41][5];
              muxOutConnector[48] = fifoOut[42][5];
              muxOutConnector[49] = fifoOut[43][5];
              muxOutConnector[50] = fifoOut[44][5];
              muxOutConnector[51] = fifoOut[45][5];
       end
       14: begin
              muxOutConnector[0] = fifoOut[1][3];
              muxOutConnector[1] = fifoOut[2][3];
              muxOutConnector[2] = fifoOut[3][3];
              muxOutConnector[3] = fifoOut[4][3];
              muxOutConnector[4] = fifoOut[5][3];
              muxOutConnector[5] = fifoOut[6][3];
              muxOutConnector[6] = fifoOut[7][3];
              muxOutConnector[7] = fifoOut[8][3];
              muxOutConnector[8] = fifoOut[9][3];
              muxOutConnector[9] = fifoOut[10][3];
              muxOutConnector[10] = fifoOut[11][3];
              muxOutConnector[11] = fifoOut[12][3];
              muxOutConnector[12] = fifoOut[13][3];
              muxOutConnector[13] = fifoOut[14][3];
              muxOutConnector[14] = fifoOut[15][3];
              muxOutConnector[15] = fifoOut[16][3];
              muxOutConnector[16] = fifoOut[45][2];
              muxOutConnector[17] = fifoOut[46][2];
              muxOutConnector[18] = fifoOut[47][2];
              muxOutConnector[19] = fifoOut[48][2];
              muxOutConnector[20] = fifoOut[49][2];
              muxOutConnector[21] = fifoOut[50][2];
              muxOutConnector[22] = fifoOut[51][2];
              muxOutConnector[23] = fifoOut[26][1];
              muxOutConnector[24] = fifoOut[27][1];
              muxOutConnector[25] = fifoOut[28][1];
              muxOutConnector[26] = fifoOut[46][6];
              muxOutConnector[27] = fifoOut[47][6];
              muxOutConnector[28] = fifoOut[48][6];
              muxOutConnector[29] = fifoOut[49][6];
              muxOutConnector[30] = fifoOut[50][6];
              muxOutConnector[31] = fifoOut[51][6];
              muxOutConnector[32] = fifoOut[26][5];
              muxOutConnector[33] = fifoOut[27][5];
              muxOutConnector[34] = fifoOut[28][5];
              muxOutConnector[35] = fifoOut[29][5];
              muxOutConnector[36] = fifoOut[30][5];
              muxOutConnector[37] = fifoOut[31][5];
              muxOutConnector[38] = fifoOut[32][5];
              muxOutConnector[39] = fifoOut[33][5];
              muxOutConnector[40] = fifoOut[34][5];
              muxOutConnector[41] = fifoOut[35][5];
              muxOutConnector[42] = fifoOut[36][5];
              muxOutConnector[43] = fifoOut[37][5];
              muxOutConnector[44] = fifoOut[38][5];
              muxOutConnector[45] = fifoOut[39][5];
              muxOutConnector[46] = fifoOut[40][5];
              muxOutConnector[47] = fifoOut[41][5];
              muxOutConnector[48] = fifoOut[42][5];
              muxOutConnector[49] = fifoOut[43][5];
              muxOutConnector[50] = fifoOut[44][5];
              muxOutConnector[51] = fifoOut[45][5];
       end
       15: begin
              muxOutConnector[0] = fifoOut[29][2];
              muxOutConnector[1] = fifoOut[30][2];
              muxOutConnector[2] = fifoOut[31][2];
              muxOutConnector[3] = fifoOut[32][2];
              muxOutConnector[4] = fifoOut[33][2];
              muxOutConnector[5] = fifoOut[34][2];
              muxOutConnector[6] = fifoOut[35][2];
              muxOutConnector[7] = fifoOut[36][2];
              muxOutConnector[8] = fifoOut[37][2];
              muxOutConnector[9] = fifoOut[38][2];
              muxOutConnector[10] = fifoOut[39][2];
              muxOutConnector[11] = fifoOut[40][2];
              muxOutConnector[12] = fifoOut[41][2];
              muxOutConnector[13] = fifoOut[42][2];
              muxOutConnector[14] = fifoOut[43][2];
              muxOutConnector[15] = fifoOut[44][2];
              muxOutConnector[16] = fifoOut[45][2];
              muxOutConnector[17] = fifoOut[46][2];
              muxOutConnector[18] = fifoOut[47][2];
              muxOutConnector[19] = fifoOut[48][2];
              muxOutConnector[20] = fifoOut[49][2];
              muxOutConnector[21] = fifoOut[50][2];
              muxOutConnector[22] = fifoOut[51][2];
              muxOutConnector[23] = fifoOut[26][1];
              muxOutConnector[24] = fifoOut[27][1];
              muxOutConnector[25] = fifoOut[28][1];
              muxOutConnector[26] = fifoOut[46][6];
              muxOutConnector[27] = fifoOut[47][6];
              muxOutConnector[28] = fifoOut[48][6];
              muxOutConnector[29] = fifoOut[49][6];
              muxOutConnector[30] = fifoOut[50][6];
              muxOutConnector[31] = fifoOut[51][6];
              muxOutConnector[32] = fifoOut[26][5];
              muxOutConnector[33] = fifoOut[27][5];
              muxOutConnector[34] = fifoOut[28][5];
              muxOutConnector[35] = fifoOut[29][5];
              muxOutConnector[36] = fifoOut[30][5];
              muxOutConnector[37] = fifoOut[31][5];
              muxOutConnector[38] = fifoOut[32][5];
              muxOutConnector[39] = fifoOut[33][5];
              muxOutConnector[40] = fifoOut[34][5];
              muxOutConnector[41] = fifoOut[35][5];
              muxOutConnector[42] = fifoOut[36][5];
              muxOutConnector[43] = fifoOut[37][5];
              muxOutConnector[44] = fifoOut[38][5];
              muxOutConnector[45] = fifoOut[39][5];
              muxOutConnector[46] = fifoOut[40][5];
              muxOutConnector[47] = fifoOut[41][5];
              muxOutConnector[48] = fifoOut[42][5];
              muxOutConnector[49] = fifoOut[43][5];
              muxOutConnector[50] = fifoOut[44][5];
              muxOutConnector[51] = fifoOut[45][5];
       end
       16: begin
              muxOutConnector[0] = fifoOut[29][2];
              muxOutConnector[1] = fifoOut[30][2];
              muxOutConnector[2] = fifoOut[31][2];
              muxOutConnector[3] = fifoOut[32][2];
              muxOutConnector[4] = fifoOut[33][2];
              muxOutConnector[5] = fifoOut[34][2];
              muxOutConnector[6] = fifoOut[35][2];
              muxOutConnector[7] = fifoOut[36][2];
              muxOutConnector[8] = fifoOut[37][2];
              muxOutConnector[9] = fifoOut[38][2];
              muxOutConnector[10] = fifoOut[39][2];
              muxOutConnector[11] = fifoOut[40][2];
              muxOutConnector[12] = fifoOut[41][2];
              muxOutConnector[13] = fifoOut[42][2];
              muxOutConnector[14] = fifoOut[43][2];
              muxOutConnector[15] = fifoOut[44][2];
              muxOutConnector[16] = fifoOut[45][2];
              muxOutConnector[17] = fifoOut[46][2];
              muxOutConnector[18] = fifoOut[47][2];
              muxOutConnector[19] = fifoOut[48][2];
              muxOutConnector[20] = fifoOut[49][2];
              muxOutConnector[21] = fifoOut[50][2];
              muxOutConnector[22] = fifoOut[51][2];
              muxOutConnector[23] = fifoOut[26][1];
              muxOutConnector[24] = fifoOut[27][1];
              muxOutConnector[25] = fifoOut[28][1];
              muxOutConnector[26] = fifoOut[46][6];
              muxOutConnector[27] = fifoOut[47][6];
              muxOutConnector[28] = fifoOut[48][6];
              muxOutConnector[29] = fifoOut[49][6];
              muxOutConnector[30] = fifoOut[50][6];
              muxOutConnector[31] = fifoOut[51][6];
              muxOutConnector[32] = fifoOut[26][5];
              muxOutConnector[33] = fifoOut[27][5];
              muxOutConnector[34] = fifoOut[28][5];
              muxOutConnector[35] = fifoOut[29][5];
              muxOutConnector[36] = fifoOut[30][5];
              muxOutConnector[37] = fifoOut[31][5];
              muxOutConnector[38] = fifoOut[32][5];
              muxOutConnector[39] = fifoOut[33][5];
              muxOutConnector[40] = fifoOut[34][5];
              muxOutConnector[41] = fifoOut[35][5];
              muxOutConnector[42] = fifoOut[36][5];
              muxOutConnector[43] = fifoOut[37][5];
              muxOutConnector[44] = fifoOut[38][5];
              muxOutConnector[45] = fifoOut[39][5];
              muxOutConnector[46] = fifoOut[40][5];
              muxOutConnector[47] = fifoOut[41][5];
              muxOutConnector[48] = fifoOut[42][5];
              muxOutConnector[49] = fifoOut[24][4];
              muxOutConnector[50] = fifoOut[25][4];
              muxOutConnector[51] = fifoOut[0][3];
       end
       17: begin
              muxOutConnector[0] = fifoOut[29][2];
              muxOutConnector[1] = fifoOut[30][2];
              muxOutConnector[2] = fifoOut[31][2];
              muxOutConnector[3] = fifoOut[32][2];
              muxOutConnector[4] = fifoOut[33][2];
              muxOutConnector[5] = fifoOut[34][2];
              muxOutConnector[6] = fifoOut[35][2];
              muxOutConnector[7] = fifoOut[36][2];
              muxOutConnector[8] = fifoOut[37][2];
              muxOutConnector[9] = fifoOut[38][2];
              muxOutConnector[10] = fifoOut[39][2];
              muxOutConnector[11] = fifoOut[40][2];
              muxOutConnector[12] = fifoOut[41][2];
              muxOutConnector[13] = fifoOut[42][2];
              muxOutConnector[14] = fifoOut[43][2];
              muxOutConnector[15] = fifoOut[44][2];
              muxOutConnector[16] = fifoOut[45][2];
              muxOutConnector[17] = fifoOut[46][2];
              muxOutConnector[18] = fifoOut[47][2];
              muxOutConnector[19] = fifoOut[48][2];
              muxOutConnector[20] = fifoOut[49][2];
              muxOutConnector[21] = fifoOut[50][2];
              muxOutConnector[22] = fifoOut[51][2];
              muxOutConnector[23] = fifoOut[26][1];
              muxOutConnector[24] = fifoOut[27][1];
              muxOutConnector[25] = fifoOut[28][1];
              muxOutConnector[26] = fifoOut[1][4];
              muxOutConnector[27] = fifoOut[2][4];
              muxOutConnector[28] = fifoOut[3][4];
              muxOutConnector[29] = fifoOut[4][4];
              muxOutConnector[30] = fifoOut[5][4];
              muxOutConnector[31] = fifoOut[6][4];
              muxOutConnector[32] = fifoOut[7][4];
              muxOutConnector[33] = fifoOut[8][4];
              muxOutConnector[34] = fifoOut[9][4];
              muxOutConnector[35] = fifoOut[10][4];
              muxOutConnector[36] = fifoOut[11][4];
              muxOutConnector[37] = fifoOut[12][4];
              muxOutConnector[38] = fifoOut[13][4];
              muxOutConnector[39] = fifoOut[14][4];
              muxOutConnector[40] = fifoOut[15][4];
              muxOutConnector[41] = fifoOut[16][4];
              muxOutConnector[42] = fifoOut[17][4];
              muxOutConnector[43] = fifoOut[18][4];
              muxOutConnector[44] = fifoOut[19][4];
              muxOutConnector[45] = fifoOut[20][4];
              muxOutConnector[46] = fifoOut[21][4];
              muxOutConnector[47] = fifoOut[22][4];
              muxOutConnector[48] = fifoOut[23][4];
              muxOutConnector[49] = fifoOut[24][4];
              muxOutConnector[50] = fifoOut[25][4];
              muxOutConnector[51] = fifoOut[0][3];
       end
       18: begin
              muxOutConnector[0] = fifoOut[29][2];
              muxOutConnector[1] = fifoOut[30][2];
              muxOutConnector[2] = fifoOut[31][2];
              muxOutConnector[3] = fifoOut[32][2];
              muxOutConnector[4] = fifoOut[33][2];
              muxOutConnector[5] = fifoOut[34][2];
              muxOutConnector[6] = fifoOut[35][2];
              muxOutConnector[7] = fifoOut[36][2];
              muxOutConnector[8] = fifoOut[37][2];
              muxOutConnector[9] = fifoOut[38][2];
              muxOutConnector[10] = fifoOut[39][2];
              muxOutConnector[11] = fifoOut[40][2];
              muxOutConnector[12] = fifoOut[41][2];
              muxOutConnector[13] = fifoOut[42][2];
              muxOutConnector[14] = fifoOut[43][2];
              muxOutConnector[15] = fifoOut[44][2];
              muxOutConnector[16] = fifoOut[45][2];
              muxOutConnector[17] = fifoOut[46][2];
              muxOutConnector[18] = fifoOut[47][2];
              muxOutConnector[19] = fifoOut[48][2];
              muxOutConnector[20] = fifoOut[49][2];
              muxOutConnector[21] = fifoOut[50][2];
              muxOutConnector[22] = fifoOut[51][2];
              muxOutConnector[23] = fifoOut[26][1];
              muxOutConnector[24] = fifoOut[27][1];
              muxOutConnector[25] = fifoOut[28][1];
              muxOutConnector[26] = fifoOut[1][4];
              muxOutConnector[27] = fifoOut[2][4];
              muxOutConnector[28] = fifoOut[3][4];
              muxOutConnector[29] = fifoOut[4][4];
              muxOutConnector[30] = fifoOut[5][4];
              muxOutConnector[31] = fifoOut[6][4];
              muxOutConnector[32] = fifoOut[7][4];
              muxOutConnector[33] = fifoOut[8][4];
              muxOutConnector[34] = fifoOut[9][4];
              muxOutConnector[35] = fifoOut[10][4];
              muxOutConnector[36] = fifoOut[11][4];
              muxOutConnector[37] = fifoOut[12][4];
              muxOutConnector[38] = fifoOut[13][4];
              muxOutConnector[39] = fifoOut[14][4];
              muxOutConnector[40] = fifoOut[15][4];
              muxOutConnector[41] = fifoOut[16][4];
              muxOutConnector[42] = fifoOut[17][4];
              muxOutConnector[43] = fifoOut[18][4];
              muxOutConnector[44] = fifoOut[19][4];
              muxOutConnector[45] = fifoOut[20][4];
              muxOutConnector[46] = fifoOut[21][4];
              muxOutConnector[47] = fifoOut[22][4];
              muxOutConnector[48] = fifoOut[23][4];
              muxOutConnector[49] = fifoOut[24][4];
              muxOutConnector[50] = fifoOut[25][4];
              muxOutConnector[51] = fifoOut[0][3];
       end
       19: begin
              muxOutConnector[0] = fifoOut[29][2];
              muxOutConnector[1] = fifoOut[30][2];
              muxOutConnector[2] = fifoOut[31][2];
              muxOutConnector[3] = fifoOut[32][2];
              muxOutConnector[4] = fifoOut[33][2];
              muxOutConnector[5] = fifoOut[34][2];
              muxOutConnector[6] = fifoOut[35][2];
              muxOutConnector[7] = fifoOut[36][2];
              muxOutConnector[8] = fifoOut[37][2];
              muxOutConnector[9] = fifoOut[38][2];
              muxOutConnector[10] = fifoOut[39][2];
              muxOutConnector[11] = fifoOut[40][2];
              muxOutConnector[12] = fifoOut[41][2];
              muxOutConnector[13] = fifoOut[42][2];
              muxOutConnector[14] = fifoOut[43][2];
              muxOutConnector[15] = fifoOut[44][2];
              muxOutConnector[16] = fifoOut[45][2];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[1][4];
              muxOutConnector[27] = fifoOut[2][4];
              muxOutConnector[28] = fifoOut[3][4];
              muxOutConnector[29] = fifoOut[4][4];
              muxOutConnector[30] = fifoOut[5][4];
              muxOutConnector[31] = fifoOut[6][4];
              muxOutConnector[32] = fifoOut[7][4];
              muxOutConnector[33] = fifoOut[8][4];
              muxOutConnector[34] = fifoOut[9][4];
              muxOutConnector[35] = fifoOut[10][4];
              muxOutConnector[36] = fifoOut[11][4];
              muxOutConnector[37] = fifoOut[12][4];
              muxOutConnector[38] = fifoOut[13][4];
              muxOutConnector[39] = fifoOut[14][4];
              muxOutConnector[40] = fifoOut[15][4];
              muxOutConnector[41] = fifoOut[16][4];
              muxOutConnector[42] = fifoOut[17][4];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
