`timescale 1ns / 1ps
module LMem1To0_511_circ0_combined_ys_yu_scripted(
        unloadMuxOut,
        unload_en,
        unloadAddress,
        muxOut,
        ly0In,
        rxIn,
        load_input_en,
        iteration_0_indicator,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
        feedback_en,
parameter w = 6; // DataWidth
parameter r = 52;
parameter r_lower = 32;
parameter c = 17;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter unloadMuxOutBits = 32;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input load_input_en;
input iteration_0_indicator;
input [ADDRESSWIDTH-1:0]unloadAddress;
input feedback_en;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output reg [unloadMuxOutBits - 1:0]unloadMuxOut;
input unload_en;
input [ADDRESSWIDTH-1:0]unloadAddress;
output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input [ r_lower * w - 1 : 0 ] rxIn; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [ADDRESSWIDTH-1:0]unloadAddress_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
wire [w-1:0]rxInConnector[r_lower-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

generate
    for (k=0;k<r_lower;k=k+1)begin:assign_input
        assign rxInConnector[k] = rxIn[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            if(feedback_en)begin
                 fifoOut[i][0] <= fifoOut[i][c-1];
            end
            else if(load_input_en)begin
                 if(i < r_lower)begin
                   fifoOut[i][0] = rxIn[i];
                 end
                 else begin
                   fifoOut[i][0] = maxVal
                 end
            end
            else begin
                 fifoOut[i][0] <= ly0InConnector[i];
            end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

assign unloadAddress_case = unload_en ? unloadAddress : READDISABLEDCASE;

always@(*)begin
    case(unloadAddress_case)
fifoOut[25][4][w-1];
              unloadMuxOut[4] = fifoOut[0][3][w-1];
              unloadMuxOut[5] = fifoOut[1][3][w-1];
              unloadMuxOut[6] = fifoOut[2][3][w-1];
              unloadMuxOut[7] = fifoOut[3][3][w-1];
              unloadMuxOut[8] = fifoOut[4][3][w-1];
              unloadMuxOut[9] = fifoOut[5][3][w-1];
              unloadMuxOut[10] = fifoOut[6][3][w-1];
              unloadMuxOut[11] = fifoOut[7][3][w-1];
              unloadMuxOut[12] = fifoOut[8][3][w-1];
              unloadMuxOut[13] = fifoOut[9][3][w-1];
              unloadMuxOut[14] = fifoOut[10][3][w-1];
              unloadMuxOut[15] = fifoOut[11][3][w-1];
              unloadMuxOut[16] = fifoOut[12][3][w-1];
              unloadMuxOut[17] = fifoOut[13][3][w-1];
              unloadMuxOut[18] = fifoOut[14][3][w-1];
              unloadMuxOut[19] = fifoOut[15][3][w-1];
              unloadMuxOut[20] = fifoOut[16][3][w-1];
              unloadMuxOut[21] = fifoOut[17][3][w-1];
              unloadMuxOut[22] = fifoOut[18][3][w-1];
              unloadMuxOut[23] = fifoOut[19][3][w-1];
              unloadMuxOut[24] = fifoOut[20][3][w-1];
              unloadMuxOut[25] = fifoOut[21][3][w-1];
              unloadMuxOut[26] = fifoOut[22][3][w-1];
              unloadMuxOut[27] = fifoOut[23][3][w-1];
              unloadMuxOut[28] = fifoOut[24][3][w-1];
              unloadMuxOut[29] = fifoOut[25][3][w-1];
              unloadMuxOut[30] = fifoOut[0][2][w-1];
              unloadMuxOut[31] = fifoOut[1][2][w-1];
       end
       1: begin
              unloadMuxOut[0] = fifoOut[2][3][w-1];
              unloadMuxOut[1] = fifoOut[3][3][w-1];
              unloadMuxOut[2] = fifoOut[4][3][w-1];
              unloadMuxOut[3] = fifoOut[5][3][w-1];
              unloadMuxOut[4] = fifoOut[6][3][w-1];
              unloadMuxOut[5] = fifoOut[7][3][w-1];
              unloadMuxOut[6] = fifoOut[8][3][w-1];
              unloadMuxOut[7] = fifoOut[9][3][w-1];
              unloadMuxOut[8] = fifoOut[10][3][w-1];
              unloadMuxOut[9] = fifoOut[11][3][w-1];
              unloadMuxOut[10] = fifoOut[12][3][w-1];
              unloadMuxOut[11] = fifoOut[13][3][w-1];
              unloadMuxOut[12] = fifoOut[14][3][w-1];
              unloadMuxOut[13] = fifoOut[15][3][w-1];
              unloadMuxOut[14] = fifoOut[16][3][w-1];
              unloadMuxOut[15] = fifoOut[17][3][w-1];
              unloadMuxOut[16] = fifoOut[18][3][w-1];
              unloadMuxOut[17] = fifoOut[19][3][w-1];
              unloadMuxOut[18] = fifoOut[20][3][w-1];
              unloadMuxOut[19] = fifoOut[21][3][w-1];
              unloadMuxOut[20] = fifoOut[22][3][w-1];
              unloadMuxOut[21] = fifoOut[23][3][w-1];
              unloadMuxOut[22] = fifoOut[24][3][w-1];
              unloadMuxOut[23] = fifoOut[25][3][w-1];
              unloadMuxOut[24] = fifoOut[0][2][w-1];
              unloadMuxOut[25] = fifoOut[1][2][w-1];
              unloadMuxOut[26] = fifoOut[2][2][w-1];
              unloadMuxOut[27] = fifoOut[3][2][w-1];
              unloadMuxOut[28] = fifoOut[4][2][w-1];
              unloadMuxOut[29] = fifoOut[5][2][w-1];
              unloadMuxOut[30] = fifoOut[6][2][w-1];
              unloadMuxOut[31] = fifoOut[7][2][w-1];
       end
       2: begin
              unloadMuxOut[0] = fifoOut[8][3][w-1];
              unloadMuxOut[1] = fifoOut[9][3][w-1];
              unloadMuxOut[2] = fifoOut[10][3][w-1];
              unloadMuxOut[3] = fifoOut[11][3][w-1];
              unloadMuxOut[4] = fifoOut[12][3][w-1];
              unloadMuxOut[5] = fifoOut[13][3][w-1];
              unloadMuxOut[6] = fifoOut[14][3][w-1];
              unloadMuxOut[7] = fifoOut[15][3][w-1];
              unloadMuxOut[8] = fifoOut[16][3][w-1];
              unloadMuxOut[9] = fifoOut[17][3][w-1];
              unloadMuxOut[10] = fifoOut[18][3][w-1];
              unloadMuxOut[11] = fifoOut[19][3][w-1];
              unloadMuxOut[12] = fifoOut[20][3][w-1];
              unloadMuxOut[13] = fifoOut[21][3][w-1];
              unloadMuxOut[14] = fifoOut[22][3][w-1];
              unloadMuxOut[15] = fifoOut[23][3][w-1];
              unloadMuxOut[16] = fifoOut[24][3][w-1];
              unloadMuxOut[17] = fifoOut[25][3][w-1];
              unloadMuxOut[18] = fifoOut[0][2][w-1];
              unloadMuxOut[19] = fifoOut[1][2][w-1];
              unloadMuxOut[20] = fifoOut[2][2][w-1];
              unloadMuxOut[21] = fifoOut[3][2][w-1];
              unloadMuxOut[22] = fifoOut[4][2][w-1];
              unloadMuxOut[23] = fifoOut[5][2][w-1];
              unloadMuxOut[24] = fifoOut[6][2][w-1];
              unloadMuxOut[25] = fifoOut[7][2][w-1];
              unloadMuxOut[26] = fifoOut[26][16][w-1];
              unloadMuxOut[27] = fifoOut[27][16][w-1];
              unloadMuxOut[28] = fifoOut[28][16][w-1];
              unloadMuxOut[29] = fifoOut[29][16][w-1];
              unloadMuxOut[30] = fifoOut[30][16][w-1];
              unloadMuxOut[31] = fifoOut[31][16][w-1];
       end
       3: begin
              unloadMuxOut[0] = fifoOut[14][3][w-1];
              unloadMuxOut[1] = fifoOut[15][3][w-1];
              unloadMuxOut[2] = fifoOut[16][3][w-1];
              unloadMuxOut[3] = fifoOut[35][0][w-1];
              unloadMuxOut[4] = fifoOut[36][0][w-1];
              unloadMuxOut[5] = fifoOut[37][0][w-1];
              unloadMuxOut[6] = fifoOut[38][0][w-1];
              unloadMuxOut[7] = fifoOut[39][0][w-1];
              unloadMuxOut[8] = fifoOut[40][0][w-1];
              unloadMuxOut[9] = fifoOut[41][0][w-1];
              unloadMuxOut[10] = fifoOut[42][0][w-1];
              unloadMuxOut[11] = fifoOut[43][0][w-1];
              unloadMuxOut[12] = fifoOut[44][0][w-1];
              unloadMuxOut[13] = fifoOut[45][0][w-1];
              unloadMuxOut[14] = fifoOut[46][0][w-1];
              unloadMuxOut[15] = fifoOut[47][0][w-1];
              unloadMuxOut[16] = fifoOut[48][0][w-1];
              unloadMuxOut[17] = fifoOut[49][0][w-1];
              unloadMuxOut[18] = fifoOut[50][0][w-1];
              unloadMuxOut[19] = fifoOut[51][0][w-1];
              unloadMuxOut[20] = fifoOut[26][16][w-1];
              unloadMuxOut[21] = fifoOut[27][16][w-1];
              unloadMuxOut[22] = fifoOut[28][16][w-1];
              unloadMuxOut[23] = fifoOut[29][16][w-1];
              unloadMuxOut[24] = fifoOut[30][16][w-1];
              unloadMuxOut[25] = fifoOut[31][16][w-1];
              unloadMuxOut[26] = fifoOut[32][16][w-1];
              unloadMuxOut[27] = fifoOut[33][16][w-1];
              unloadMuxOut[28] = fifoOut[34][16][w-1];
              unloadMuxOut[29] = fifoOut[35][16][w-1];
              unloadMuxOut[30] = fifoOut[36][16][w-1];
              unloadMuxOut[31] = fifoOut[37][16][w-1];
       end
       4: begin
              unloadMuxOut[0] = fifoOut[38][0][w-1];
              unloadMuxOut[1] = fifoOut[39][0][w-1];
              unloadMuxOut[2] = fifoOut[40][0][w-1];
              unloadMuxOut[3] = fifoOut[41][0][w-1];
              unloadMuxOut[4] = fifoOut[42][0][w-1];
              unloadMuxOut[5] = fifoOut[43][0][w-1];
              unloadMuxOut[6] = fifoOut[44][0][w-1];
              unloadMuxOut[7] = fifoOut[45][0][w-1];
              unloadMuxOut[8] = fifoOut[46][0][w-1];
              unloadMuxOut[9] = fifoOut[47][0][w-1];
              unloadMuxOut[10] = fifoOut[48][0][w-1];
              unloadMuxOut[11] = fifoOut[49][0][w-1];
              unloadMuxOut[12] = fifoOut[50][0][w-1];
              unloadMuxOut[13] = fifoOut[51][0][w-1];
              unloadMuxOut[14] = fifoOut[26][16][w-1];
              unloadMuxOut[15] = fifoOut[27][16][w-1];
              unloadMuxOut[16] = fifoOut[28][16][w-1];
              unloadMuxOut[17] = fifoOut[29][16][w-1];
              unloadMuxOut[18] = fifoOut[30][16][w-1];
              unloadMuxOut[19] = fifoOut[31][16][w-1];
              unloadMuxOut[20] = fifoOut[32][16][w-1];
              unloadMuxOut[21] = fifoOut[33][16][w-1];
              unloadMuxOut[22] = fifoOut[34][16][w-1];
              unloadMuxOut[23] = fifoOut[35][16][w-1];
              unloadMuxOut[24] = fifoOut[36][16][w-1];
              unloadMuxOut[25] = fifoOut[37][16][w-1];
              unloadMuxOut[26] = fifoOut[38][16][w-1];
              unloadMuxOut[27] = fifoOut[39][16][w-1];
              unloadMuxOut[28] = fifoOut[40][16][w-1];
              unloadMuxOut[29] = fifoOut[41][16][w-1];
              unloadMuxOut[30] = fifoOut[42][16][w-1];
              unloadMuxOut[31] = fifoOut[43][16][w-1];
       end
       5: begin
              unloadMuxOut[0] = fifoOut[44][0][w-1];
              unloadMuxOut[1] = fifoOut[45][0][w-1];
              unloadMuxOut[2] = fifoOut[46][0][w-1];
              unloadMuxOut[3] = fifoOut[47][0][w-1];
              unloadMuxOut[4] = fifoOut[48][0][w-1];
              unloadMuxOut[5] = fifoOut[49][0][w-1];
              unloadMuxOut[6] = fifoOut[50][0][w-1];
              unloadMuxOut[7] = fifoOut[51][0][w-1];
              unloadMuxOut[8] = fifoOut[26][16][w-1];
              unloadMuxOut[9] = fifoOut[27][16][w-1];
              unloadMuxOut[10] = fifoOut[28][16][w-1];
              unloadMuxOut[11] = fifoOut[29][16][w-1];
              unloadMuxOut[12] = fifoOut[30][16][w-1];
              unloadMuxOut[13] = fifoOut[31][16][w-1];
              unloadMuxOut[14] = fifoOut[32][16][w-1];
              unloadMuxOut[15] = fifoOut[33][16][w-1];
              unloadMuxOut[16] = fifoOut[34][16][w-1];
              unloadMuxOut[17] = fifoOut[35][16][w-1];
              unloadMuxOut[18] = fifoOut[36][16][w-1];
              unloadMuxOut[19] = fifoOut[37][16][w-1];
              unloadMuxOut[20] = fifoOut[38][16][w-1];
              unloadMuxOut[21] = fifoOut[39][16][w-1];
              unloadMuxOut[22] = fifoOut[40][16][w-1];
              unloadMuxOut[23] = fifoOut[41][16][w-1];
              unloadMuxOut[24] = fifoOut[42][16][w-1];
              unloadMuxOut[25] = fifoOut[43][16][w-1];
              unloadMuxOut[26] = fifoOut[44][16][w-1];
              unloadMuxOut[27] = fifoOut[45][16][w-1];
              unloadMuxOut[28] = fifoOut[46][16][w-1];
              unloadMuxOut[29] = fifoOut[47][16][w-1];
              unloadMuxOut[30] = fifoOut[48][16][w-1];
              unloadMuxOut[31] = fifoOut[49][16][w-1];
       end
       6: begin
              unloadMuxOut[0] = fifoOut[50][0][w-1];
              unloadMuxOut[1] = fifoOut[51][0][w-1];
              unloadMuxOut[2] = fifoOut[26][16][w-1];
              unloadMuxOut[3] = fifoOut[27][16][w-1];
              unloadMuxOut[4] = fifoOut[28][16][w-1];
              unloadMuxOut[5] = fifoOut[29][16][w-1];
              unloadMuxOut[6] = fifoOut[30][16][w-1];
              unloadMuxOut[7] = fifoOut[31][16][w-1];
              unloadMuxOut[8] = fifoOut[32][16][w-1];
              unloadMuxOut[9] = fifoOut[33][16][w-1];
              unloadMuxOut[10] = fifoOut[34][16][w-1];
              unloadMuxOut[11] = fifoOut[35][16][w-1];
              unloadMuxOut[12] = fifoOut[36][16][w-1];
              unloadMuxOut[13] = fifoOut[37][16][w-1];
              unloadMuxOut[14] = fifoOut[38][16][w-1];
              unloadMuxOut[15] = fifoOut[39][16][w-1];
              unloadMuxOut[16] = fifoOut[40][16][w-1];
              unloadMuxOut[17] = fifoOut[41][16][w-1];
              unloadMuxOut[18] = fifoOut[42][16][w-1];
              unloadMuxOut[19] = fifoOut[43][16][w-1];
              unloadMuxOut[20] = fifoOut[44][16][w-1];
              unloadMuxOut[21] = fifoOut[45][16][w-1];
              unloadMuxOut[22] = fifoOut[46][16][w-1];
              unloadMuxOut[23] = fifoOut[47][16][w-1];
              unloadMuxOut[24] = fifoOut[48][16][w-1];
              unloadMuxOut[25] = fifoOut[49][16][w-1];
              unloadMuxOut[26] = fifoOut[50][16][w-1];
              unloadMuxOut[27] = fifoOut[51][16][w-1];
              unloadMuxOut[28] = fifoOut[26][15][w-1];
              unloadMuxOut[29] = fifoOut[27][15][w-1];
              unloadMuxOut[30] = fifoOut[28][15][w-1];
              unloadMuxOut[31] = fifoOut[29][15][w-1];
       end
       7: begin
              unloadMuxOut[0] = fifoOut[30][16][w-1];
              unloadMuxOut[1] = fifoOut[31][16][w-1];
              unloadMuxOut[2] = fifoOut[32][16][w-1];
              unloadMuxOut[3] = fifoOut[33][16][w-1];
              unloadMuxOut[4] = fifoOut[34][16][w-1];
              unloadMuxOut[5] = fifoOut[35][16][w-1];
              unloadMuxOut[6] = fifoOut[36][16][w-1];
              unloadMuxOut[7] = fifoOut[37][16][w-1];
              unloadMuxOut[8] = fifoOut[38][16][w-1];
              unloadMuxOut[9] = fifoOut[39][16][w-1];
              unloadMuxOut[10] = fifoOut[40][16][w-1];
              unloadMuxOut[11] = fifoOut[41][16][w-1];
              unloadMuxOut[12] = fifoOut[42][16][w-1];
              unloadMuxOut[13] = fifoOut[43][16][w-1];
              unloadMuxOut[14] = fifoOut[44][16][w-1];
              unloadMuxOut[15] = fifoOut[45][16][w-1];
              unloadMuxOut[16] = fifoOut[46][16][w-1];
              unloadMuxOut[17] = fifoOut[47][16][w-1];
              unloadMuxOut[18] = fifoOut[48][16][w-1];
              unloadMuxOut[19] = fifoOut[49][16][w-1];
              unloadMuxOut[20] = fifoOut[50][16][w-1];
              unloadMuxOut[21] = fifoOut[51][16][w-1];
              unloadMuxOut[22] = fifoOut[26][15][w-1];
              unloadMuxOut[23] = fifoOut[27][15][w-1];
              unloadMuxOut[24] = fifoOut[28][15][w-1];
              unloadMuxOut[25] = fifoOut[29][15][w-1];
              unloadMuxOut[26] = fifoOut[30][15][w-1];
              unloadMuxOut[27] = fifoOut[31][15][w-1];
              unloadMuxOut[28] = fifoOut[32][15][w-1];
              unloadMuxOut[29] = fifoOut[33][15][w-1];
              unloadMuxOut[30] = fifoOut[34][15][w-1];
              unloadMuxOut[31] = fifoOut[35][15][w-1];
       end
       8: begin
              unloadMuxOut[0] = fifoOut[36][16][w-1];
              unloadMuxOut[1] = fifoOut[37][16][w-1];
              unloadMuxOut[2] = fifoOut[38][16][w-1];
              unloadMuxOut[3] = fifoOut[39][16][w-1];
              unloadMuxOut[4] = fifoOut[40][16][w-1];
              unloadMuxOut[5] = fifoOut[41][16][w-1];
              unloadMuxOut[6] = fifoOut[42][16][w-1];
              unloadMuxOut[7] = fifoOut[43][16][w-1];
              unloadMuxOut[8] = fifoOut[44][16][w-1];
              unloadMuxOut[9] = fifoOut[45][16][w-1];
              unloadMuxOut[10] = fifoOut[46][16][w-1];
              unloadMuxOut[11] = fifoOut[47][16][w-1];
              unloadMuxOut[12] = fifoOut[48][16][w-1];
              unloadMuxOut[13] = fifoOut[49][16][w-1];
              unloadMuxOut[14] = fifoOut[50][16][w-1];
              unloadMuxOut[15] = fifoOut[51][16][w-1];
              unloadMuxOut[16] = fifoOut[26][15][w-1];
              unloadMuxOut[17] = fifoOut[27][15][w-1];
              unloadMuxOut[18] = fifoOut[28][15][w-1];
              unloadMuxOut[19] = fifoOut[29][15][w-1];
              unloadMuxOut[20] = fifoOut[30][15][w-1];
              unloadMuxOut[21] = fifoOut[31][15][w-1];
              unloadMuxOut[22] = fifoOut[32][15][w-1];
              unloadMuxOut[23] = fifoOut[33][15][w-1];
              unloadMuxOut[24] = fifoOut[34][15][w-1];
              unloadMuxOut[25] = fifoOut[35][15][w-1];
              unloadMuxOut[26] = fifoOut[36][15][w-1];
              unloadMuxOut[27] = fifoOut[37][15][w-1];
              unloadMuxOut[28] = fifoOut[38][15][w-1];
              unloadMuxOut[29] = fifoOut[39][15][w-1];
              unloadMuxOut[30] = fifoOut[40][15][w-1];
              unloadMuxOut[31] = fifoOut[41][15][w-1];
       end
       9: begin
              unloadMuxOut[0] = fifoOut[42][16][w-1];
              unloadMuxOut[1] = fifoOut[43][16][w-1];
              unloadMuxOut[2] = fifoOut[44][16][w-1];
              unloadMuxOut[3] = fifoOut[45][16][w-1];
              unloadMuxOut[4] = fifoOut[46][16][w-1];
              unloadMuxOut[5] = fifoOut[47][16][w-1];
              unloadMuxOut[6] = fifoOut[48][16][w-1];
              unloadMuxOut[7] = fifoOut[49][16][w-1];
              unloadMuxOut[8] = fifoOut[50][16][w-1];
              unloadMuxOut[9] = fifoOut[51][16][w-1];
              unloadMuxOut[10] = fifoOut[26][15][w-1];
              unloadMuxOut[11] = fifoOut[27][15][w-1];
              unloadMuxOut[12] = fifoOut[28][15][w-1];
              unloadMuxOut[13] = fifoOut[29][15][w-1];
              unloadMuxOut[14] = fifoOut[30][15][w-1];
              unloadMuxOut[15] = fifoOut[31][15][w-1];
              unloadMuxOut[16] = fifoOut[32][15][w-1];
              unloadMuxOut[17] = fifoOut[33][15][w-1];
              unloadMuxOut[18] = fifoOut[34][15][w-1];
              unloadMuxOut[19] = fifoOut[35][15][w-1];
              unloadMuxOut[20] = fifoOut[36][15][w-1];
              unloadMuxOut[21] = fifoOut[37][15][w-1];
              unloadMuxOut[22] = fifoOut[38][15][w-1];
              unloadMuxOut[23] = fifoOut[39][15][w-1];
              unloadMuxOut[24] = fifoOut[40][15][w-1];
              unloadMuxOut[25] = fifoOut[41][15][w-1];
              unloadMuxOut[26] = fifoOut[42][15][w-1];
              unloadMuxOut[27] = fifoOut[43][15][w-1];
              unloadMuxOut[28] = fifoOut[44][15][w-1];
              unloadMuxOut[29] = fifoOut[45][15][w-1];
              unloadMuxOut[30] = fifoOut[46][15][w-1];
              unloadMuxOut[31] = fifoOut[47][15][w-1];
       end
       10: begin
              unloadMuxOut[0] = fifoOut[48][16][w-1];
              unloadMuxOut[1] = fifoOut[49][16][w-1];
              unloadMuxOut[2] = fifoOut[50][16][w-1];
              unloadMuxOut[3] = fifoOut[51][16][w-1];
              unloadMuxOut[4] = fifoOut[26][15][w-1];
              unloadMuxOut[5] = fifoOut[27][15][w-1];
              unloadMuxOut[6] = fifoOut[28][15][w-1];
              unloadMuxOut[7] = fifoOut[29][15][w-1];
              unloadMuxOut[8] = fifoOut[30][15][w-1];
              unloadMuxOut[9] = fifoOut[31][15][w-1];
              unloadMuxOut[10] = fifoOut[32][15][w-1];
              unloadMuxOut[11] = fifoOut[33][15][w-1];
              unloadMuxOut[12] = fifoOut[34][15][w-1];
              unloadMuxOut[13] = fifoOut[35][15][w-1];
              unloadMuxOut[14] = fifoOut[36][15][w-1];
              unloadMuxOut[15] = fifoOut[37][15][w-1];
              unloadMuxOut[16] = fifoOut[38][15][w-1];
              unloadMuxOut[17] = fifoOut[39][15][w-1];
              unloadMuxOut[18] = fifoOut[40][15][w-1];
              unloadMuxOut[19] = fifoOut[41][15][w-1];
              unloadMuxOut[20] = fifoOut[42][15][w-1];
              unloadMuxOut[21] = fifoOut[43][15][w-1];
              unloadMuxOut[22] = fifoOut[44][15][w-1];
              unloadMuxOut[23] = fifoOut[45][15][w-1];
              unloadMuxOut[24] = fifoOut[46][15][w-1];
              unloadMuxOut[25] = fifoOut[47][15][w-1];
              unloadMuxOut[26] = fifoOut[48][15][w-1];
              unloadMuxOut[27] = fifoOut[49][15][w-1];
              unloadMuxOut[28] = fifoOut[50][15][w-1];
              unloadMuxOut[29] = fifoOut[51][15][w-1];
              unloadMuxOut[30] = fifoOut[26][14][w-1];
              unloadMuxOut[31] = fifoOut[27][14][w-1];
       end
       11: begin
              unloadMuxOut[0] = fifoOut[28][15][w-1];
              unloadMuxOut[1] = fifoOut[29][15][w-1];
              unloadMuxOut[2] = fifoOut[30][15][w-1];
              unloadMuxOut[3] = fifoOut[31][15][w-1];
              unloadMuxOut[4] = fifoOut[32][15][w-1];
              unloadMuxOut[5] = fifoOut[33][15][w-1];
              unloadMuxOut[6] = fifoOut[34][15][w-1];
              unloadMuxOut[7] = fifoOut[35][15][w-1];
              unloadMuxOut[8] = fifoOut[36][15][w-1];
              unloadMuxOut[9] = fifoOut[37][15][w-1];
              unloadMuxOut[10] = fifoOut[38][15][w-1];
              unloadMuxOut[11] = fifoOut[39][15][w-1];
              unloadMuxOut[12] = fifoOut[40][15][w-1];
              unloadMuxOut[13] = fifoOut[41][15][w-1];
              unloadMuxOut[14] = fifoOut[42][15][w-1];
              unloadMuxOut[15] = fifoOut[43][15][w-1];
              unloadMuxOut[16] = fifoOut[44][15][w-1];
              unloadMuxOut[17] = fifoOut[45][15][w-1];
              unloadMuxOut[18] = fifoOut[46][15][w-1];
              unloadMuxOut[19] = fifoOut[47][15][w-1];
              unloadMuxOut[20] = fifoOut[48][15][w-1];
              unloadMuxOut[21] = fifoOut[49][15][w-1];
              unloadMuxOut[22] = fifoOut[50][15][w-1];
              unloadMuxOut[23] = fifoOut[51][15][w-1];
              unloadMuxOut[24] = fifoOut[26][14][w-1];
              unloadMuxOut[25] = fifoOut[27][14][w-1];
              unloadMuxOut[26] = fifoOut[28][14][w-1];
              unloadMuxOut[27] = fifoOut[29][14][w-1];
              unloadMuxOut[28] = fifoOut[30][14][w-1];
              unloadMuxOut[29] = fifoOut[31][14][w-1];
              unloadMuxOut[30] = fifoOut[32][14][w-1];
              unloadMuxOut[31] = fifoOut[33][14][w-1];
       end
       12: begin
              unloadMuxOut[0] = fifoOut[34][15][w-1];
              unloadMuxOut[1] = fifoOut[35][15][w-1];
              unloadMuxOut[2] = fifoOut[36][15][w-1];
              unloadMuxOut[3] = fifoOut[37][15][w-1];
              unloadMuxOut[4] = fifoOut[38][15][w-1];
              unloadMuxOut[5] = fifoOut[39][15][w-1];
              unloadMuxOut[6] = fifoOut[40][15][w-1];
              unloadMuxOut[7] = fifoOut[41][15][w-1];
              unloadMuxOut[8] = fifoOut[42][15][w-1];
              unloadMuxOut[9] = fifoOut[43][15][w-1];
              unloadMuxOut[10] = fifoOut[44][15][w-1];
              unloadMuxOut[11] = fifoOut[45][15][w-1];
              unloadMuxOut[12] = fifoOut[46][15][w-1];
              unloadMuxOut[13] = fifoOut[47][15][w-1];
              unloadMuxOut[14] = fifoOut[48][15][w-1];
              unloadMuxOut[15] = fifoOut[49][15][w-1];
              unloadMuxOut[16] = fifoOut[50][15][w-1];
              unloadMuxOut[17] = fifoOut[51][15][w-1];
              unloadMuxOut[18] = fifoOut[26][14][w-1];
              unloadMuxOut[19] = fifoOut[27][14][w-1];
              unloadMuxOut[20] = fifoOut[28][14][w-1];
              unloadMuxOut[21] = fifoOut[29][14][w-1];
              unloadMuxOut[22] = fifoOut[30][14][w-1];
              unloadMuxOut[23] = fifoOut[31][14][w-1];
              unloadMuxOut[24] = fifoOut[32][14][w-1];
              unloadMuxOut[25] = fifoOut[33][14][w-1];
              unloadMuxOut[26] = fifoOut[34][14][w-1];
              unloadMuxOut[27] = fifoOut[35][14][w-1];
              unloadMuxOut[28] = fifoOut[36][14][w-1];
              unloadMuxOut[29] = fifoOut[37][14][w-1];
              unloadMuxOut[30] = fifoOut[38][14][w-1];
              unloadMuxOut[31] = fifoOut[39][14][w-1];
       end
       13: begin
              unloadMuxOut[0] = fifoOut[40][15][w-1];
              unloadMuxOut[1] = fifoOut[41][15][w-1];
              unloadMuxOut[2] = fifoOut[42][15][w-1];
              unloadMuxOut[3] = fifoOut[43][15][w-1];
              unloadMuxOut[4] = fifoOut[44][15][w-1];
              unloadMuxOut[5] = fifoOut[45][15][w-1];
              unloadMuxOut[6] = fifoOut[46][15][w-1];
              unloadMuxOut[7] = fifoOut[47][15][w-1];
              unloadMuxOut[8] = fifoOut[48][15][w-1];
              unloadMuxOut[9] = fifoOut[49][15][w-1];
              unloadMuxOut[10] = fifoOut[50][15][w-1];
              unloadMuxOut[11] = fifoOut[51][15][w-1];
              unloadMuxOut[12] = fifoOut[26][14][w-1];
              unloadMuxOut[13] = fifoOut[27][14][w-1];
              unloadMuxOut[14] = fifoOut[28][14][w-1];
              unloadMuxOut[15] = fifoOut[29][14][w-1];
              unloadMuxOut[16] = fifoOut[30][14][w-1];
              unloadMuxOut[17] = fifoOut[31][14][w-1];
              unloadMuxOut[18] = fifoOut[32][14][w-1];
              unloadMuxOut[19] = fifoOut[33][14][w-1];
              unloadMuxOut[20] = fifoOut[34][14][w-1];
              unloadMuxOut[21] = fifoOut[35][14][w-1];
              unloadMuxOut[22] = fifoOut[36][14][w-1];
              unloadMuxOut[23] = fifoOut[37][14][w-1];
              unloadMuxOut[24] = fifoOut[38][14][w-1];
              unloadMuxOut[25] = fifoOut[39][14][w-1];
              unloadMuxOut[26] = fifoOut[40][14][w-1];
              unloadMuxOut[27] = fifoOut[41][14][w-1];
              unloadMuxOut[28] = fifoOut[42][14][w-1];
              unloadMuxOut[29] = fifoOut[43][14][w-1];
              unloadMuxOut[30] = fifoOut[44][14][w-1];
              unloadMuxOut[31] = fifoOut[45][14][w-1];
       end
       14: begin
              unloadMuxOut[0] = fifoOut[46][15][w-1];
              unloadMuxOut[1] = fifoOut[47][15][w-1];
              unloadMuxOut[2] = fifoOut[48][15][w-1];
              unloadMuxOut[3] = fifoOut[49][15][w-1];
              unloadMuxOut[4] = fifoOut[50][15][w-1];
              unloadMuxOut[5] = fifoOut[51][15][w-1];
              unloadMuxOut[6] = fifoOut[26][14][w-1];
              unloadMuxOut[7] = fifoOut[27][14][w-1];
              unloadMuxOut[8] = fifoOut[28][14][w-1];
              unloadMuxOut[9] = fifoOut[29][14][w-1];
              unloadMuxOut[10] = fifoOut[30][14][w-1];
              unloadMuxOut[11] = fifoOut[31][14][w-1];
              unloadMuxOut[12] = fifoOut[32][14][w-1];
              unloadMuxOut[13] = fifoOut[33][14][w-1];
              unloadMuxOut[14] = fifoOut[34][14][w-1];
              unloadMuxOut[15] = fifoOut[35][14][w-1];
              unloadMuxOut[16] = fifoOut[36][14][w-1];
              unloadMuxOut[17] = fifoOut[37][14][w-1];
              unloadMuxOut[18] = fifoOut[38][14][w-1];
              unloadMuxOut[19] = fifoOut[39][14][w-1];
              unloadMuxOut[20] = fifoOut[40][14][w-1];
              unloadMuxOut[21] = fifoOut[41][14][w-1];
              unloadMuxOut[22] = fifoOut[42][14][w-1];
              unloadMuxOut[23] = fifoOut[8][2][w-1];
              unloadMuxOut[24] = fifoOut[9][2][w-1];
              unloadMuxOut[25] = fifoOut[10][2][w-1];
              unloadMuxOut[26] = fifoOut[11][2][w-1];
              unloadMuxOut[27] = fifoOut[12][2][w-1];
              unloadMuxOut[28] = fifoOut[13][2][w-1];
              unloadMuxOut[29] = fifoOut[14][2][w-1];
              unloadMuxOut[30] = fifoOut[15][2][w-1];
              unloadMuxOut[31] = fifoOut[16][2][w-1];
       end
       15: begin
              unloadMuxOut[0] = fifoOut[17][3][w-1];
              unloadMuxOut[1] = fifoOut[18][3][w-1];
              unloadMuxOut[2] = fifoOut[19][3][w-1];
              unloadMuxOut[3] = fifoOut[20][3][w-1];
              unloadMuxOut[4] = fifoOut[21][3][w-1];
              unloadMuxOut[5] = fifoOut[22][3][w-1];
              unloadMuxOut[6] = fifoOut[23][3][w-1];
              unloadMuxOut[7] = fifoOut[24][3][w-1];
              unloadMuxOut[8] = fifoOut[25][3][w-1];
              unloadMuxOut[9] = fifoOut[0][2][w-1];
              unloadMuxOut[10] = fifoOut[1][2][w-1];
              unloadMuxOut[11] = fifoOut[2][2][w-1];
              unloadMuxOut[12] = fifoOut[3][2][w-1];
              unloadMuxOut[13] = fifoOut[4][2][w-1];
              unloadMuxOut[14] = fifoOut[5][2][w-1];
              unloadMuxOut[15] = fifoOut[6][2][w-1];
              unloadMuxOut[16] = fifoOut[7][2][w-1];
              unloadMuxOut[17] = fifoOut[8][2][w-1];
              unloadMuxOut[18] = fifoOut[9][2][w-1];
              unloadMuxOut[19] = fifoOut[10][2][w-1];
              unloadMuxOut[20] = fifoOut[11][2][w-1];
              unloadMuxOut[21] = fifoOut[12][2][w-1];
              unloadMuxOut[22] = fifoOut[13][2][w-1];
              unloadMuxOut[23] = fifoOut[14][2][w-1];
              unloadMuxOut[24] = fifoOut[15][2][w-1];
              unloadMuxOut[25] = fifoOut[16][2][w-1];
              unloadMuxOut[26] = fifoOut[17][2][w-1];
              unloadMuxOut[27] = fifoOut[18][2][w-1];
              unloadMuxOut[28] = fifoOut[19][2][w-1];
              unloadMuxOut[29] = fifoOut[20][2][w-1];
              unloadMuxOut[30] = fifoOut[21][2][w-1];
              unloadMuxOut[31] = 1'b0;
       end
       16: begin
              unloadMuxOut[0] = 1'b0;
              unloadMuxOut[1] = 1'b0;
              unloadMuxOut[2] = 1'b0;
              unloadMuxOut[3] = 1'b0;
              unloadMuxOut[4] = 1'b0;
              unloadMuxOut[5] = 1'b0;
              unloadMuxOut[6] = 1'b0;
              unloadMuxOut[7] = 1'b0;
              unloadMuxOut[8] = 1'b0;
              unloadMuxOut[9] = 1'b0;
              unloadMuxOut[10] = 1'b0;
              unloadMuxOut[11] = 1'b0;
              unloadMuxOut[12] = 1'b0;
              unloadMuxOut[13] = 1'b0;
              unloadMuxOut[14] = 1'b0;
              unloadMuxOut[15] = 1'b0;
              unloadMuxOut[16] = 1'b0;
              unloadMuxOut[17] = 1'b0;
              unloadMuxOut[18] = 1'b0;
              unloadMuxOut[19] = 1'b0;
              unloadMuxOut[20] = 1'b0;
              unloadMuxOut[21] = 1'b0;
              unloadMuxOut[22] = 1'b0;
              unloadMuxOut[23] = 1'b0;
              unloadMuxOut[24] = 1'b0;
              unloadMuxOut[25] = 1'b0;
              unloadMuxOut[26] = 1'b0;
              unloadMuxOut[27] = 1'b0;
              unloadMuxOut[28] = 1'b0;
              unloadMuxOut[29] = 1'b0;
              unloadMuxOut[30] = 1'b0;
              unloadMuxOut[31] = 1'b0;
       end
       default: begin
             for(i=0;i<unloadMuxOutBits;i=i+1)begin
              unloadMuxOut[i] = 0; 
             end
       end
    endcase //unload case end
    case(iteration_0_indicator)
       0: begin
         case(rd_address_case)
         0: begin
              muxOutCo        unloadMuxOut[i] = 0;
             end
       end
    endcase
    case(iteration_0_indicator)
       0: begin
         case(rd_address_case)
         0: begin
fifoOut[25][4];
              muxOutConnector[4] = fifoOut[0][3];
              muxOutConnector[5] = fifoOut[1][3];
              muxOutConnector[6] = fifoOut[2][3];
              muxOutConnector[7] = fifoOut[3][3];
              muxOutConnector[8] = fifoOut[4][3];
              muxOutConnector[9] = fifoOut[5][3];
              muxOutConnector[10] = fifoOut[6][3];
              muxOutConnector[11] = fifoOut[7][3];
              muxOutConnector[12] = fifoOut[8][3];
              muxOutConnector[13] = fifoOut[9][3];
              muxOutConnector[14] = fifoOut[10][3];
              muxOutConnector[15] = fifoOut[11][3];
              muxOutConnector[16] = fifoOut[12][3];
              muxOutConnector[17] = fifoOut[13][3];
              muxOutConnector[18] = fifoOut[14][3];
              muxOutConnector[19] = fifoOut[15][3];
              muxOutConnector[20] = fifoOut[16][3];
              muxOutConnector[21] = fifoOut[17][3];
              muxOutConnector[22] = fifoOut[18][3];
              muxOutConnector[23] = fifoOut[19][3];
              muxOutConnector[24] = fifoOut[20][3];
              muxOutConnector[25] = fifoOut[21][3];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[35][11];
              muxOutConnector[28] = fifoOut[36][11];
              muxOutConnector[29] = fifoOut[37][11];
              muxOutConnector[30] = fifoOut[38][11];
              muxOutConnector[31] = fifoOut[39][11];
              muxOutConnector[32] = fifoOut[40][11];
              muxOutConnector[33] = fifoOut[41][11];
              muxOutConnector[34] = fifoOut[42][11];
              muxOutConnector[35] = fifoOut[43][11];
              muxOutConnector[36] = fifoOut[44][11];
              muxOutConnector[37] = fifoOut[45][11];
              muxOutConnector[38] = fifoOut[46][11];
              muxOutConnector[39] = fifoOut[47][11];
              muxOutConnector[40] = fifoOut[48][11];
              muxOutConnector[41] = fifoOut[49][11];
              muxOutConnector[42] = fifoOut[50][11];
              muxOutConnector[43] = fifoOut[51][11];
              muxOutConnector[44] = fifoOut[26][10];
              muxOutConnector[45] = fifoOut[27][10];
              muxOutConnector[46] = fifoOut[28][10];
              muxOutConnector[47] = fifoOut[29][10];
              muxOutConnector[48] = fifoOut[30][10];
              muxOutConnector[49] = fifoOut[31][10];
              muxOutConnector[50] = fifoOut[32][10];
              muxOutConnector[51] = fifoOut[33][10];
         end
         1: begin
              muxOutConnector[0] = fifoOut[22][4];
              muxOutConnector[1] = fifoOut[23][4];
              muxOutConnector[2] = fifoOut[24][4];
              muxOutConnector[3] = fifoOut[25][4];
              muxOutConnector[4] = fifoOut[0][3];
              muxOutConnector[5] = fifoOut[1][3];
              muxOutConnector[6] = fifoOut[2][3];
              muxOutConnector[7] = fifoOut[3][3];
              muxOutConnector[8] = fifoOut[4][3];
              muxOutConnector[9] = fifoOut[5][3];
              muxOutConnector[10] = fifoOut[6][3];
              muxOutConnector[11] = fifoOut[7][3];
              muxOutConnector[12] = fifoOut[8][3];
              muxOutConnector[13] = fifoOut[9][3];
              muxOutConnector[14] = fifoOut[10][3];
              muxOutConnector[15] = fifoOut[11][3];
              muxOutConnector[16] = fifoOut[12][3];
              muxOutConnector[17] = fifoOut[13][3];
              muxOutConnector[18] = fifoOut[14][3];
              muxOutConnector[19] = fifoOut[15][3];
              muxOutConnector[20] = fifoOut[16][3];
              muxOutConnector[21] = fifoOut[17][3];
              muxOutConnector[22] = fifoOut[18][3];
              muxOutConnector[23] = fifoOut[19][3];
              muxOutConnector[24] = fifoOut[20][3];
              muxOutConnector[25] = fifoOut[21][3];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[35][11];
              muxOutConnector[28] = fifoOut[36][11];
              muxOutConnector[29] = fifoOut[37][11];
              muxOutConnector[30] = fifoOut[38][11];
              muxOutConnector[31] = fifoOut[39][11];
              muxOutConnector[32] = fifoOut[40][11];
              muxOutConnector[33] = fifoOut[41][11];
              muxOutConnector[34] = fifoOut[42][11];
              muxOutConnector[35] = fifoOut[43][11];
              muxOutConnector[36] = fifoOut[44][11];
              muxOutConnector[37] = fifoOut[45][11];
              muxOutConnector[38] = fifoOut[46][11];
              muxOutConnector[39] = fifoOut[47][11];
              muxOutConnector[40] = fifoOut[48][11];
              muxOutConnector[41] = fifoOut[49][11];
              muxOutConnector[42] = fifoOut[50][11];
              muxOutConnector[43] = fifoOut[51][11];
              muxOutConnector[44] = fifoOut[26][10];
              muxOutConnector[45] = fifoOut[27][10];
              muxOutConnector[46] = fifoOut[28][10];
              muxOutConnector[47] = fifoOut[29][10];
              muxOutConnector[48] = fifoOut[30][10];
              muxOutConnector[49] = fifoOut[31][10];
              muxOutConnector[50] = fifoOut[32][10];
              muxOutConnector[51] = fifoOut[33][10];
         end
         2: begin
              muxOutConnector[0] = fifoOut[22][4];
              muxOutConnector[1] = fifoOut[23][4];
              muxOutConnector[2] = fifoOut[24][4];
              muxOutConnector[3] = fifoOut[25][4];
              muxOutConnector[4] = fifoOut[0][3];
              muxOutConnector[5] = fifoOut[1][3];
              muxOutConnector[6] = fifoOut[2][3];
              muxOutConnector[7] = fifoOut[3][3];
              muxOutConnector[8] = fifoOut[4][3];
              muxOutConnector[9] = fifoOut[5][3];
              muxOutConnector[10] = fifoOut[6][3];
              muxOutConnector[11] = fifoOut[7][3];
              muxOutConnector[12] = fifoOut[8][3];
              muxOutConnector[13] = fifoOut[9][3];
              muxOutConnector[14] = fifoOut[10][3];
              muxOutConnector[15] = fifoOut[11][3];
              muxOutConnector[16] = fifoOut[12][3];
              muxOutConnector[17] = fifoOut[13][3];
              muxOutConnector[18] = fifoOut[14][3];
              muxOutConnector[19] = fifoOut[15][3];
              muxOutConnector[20] = fifoOut[16][3];
              muxOutConnector[21] = fifoOut[17][3];
              muxOutConnector[22] = fifoOut[18][3];
              muxOutConnector[23] = fifoOut[19][3];
              muxOutConnector[24] = fifoOut[20][3];
              muxOutConnector[25] = fifoOut[21][3];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[17][16];
              muxOutConnector[45] = fifoOut[18][16];
              muxOutConnector[46] = fifoOut[19][16];
              muxOutConnector[47] = fifoOut[20][16];
              muxOutConnector[48] = fifoOut[21][16];
              muxOutConnector[49] = fifoOut[22][16];
              muxOutConnector[50] = fifoOut[23][16];
              muxOutConnector[51] = fifoOut[24][16];
         end
         3: begin
              muxOutConnector[0] = fifoOut[22][4];
              muxOutConnector[1] = fifoOut[23][4];
              muxOutConnector[2] = fifoOut[24][4];
              muxOutConnector[3] = fifoOut[25][4];
              muxOutConnector[4] = fifoOut[0][3];
              muxOutConnector[5] = fifoOut[1][3];
              muxOutConnector[6] = fifoOut[2][3];
              muxOutConnector[7] = fifoOut[3][3];
              muxOutConnector[8] = fifoOut[4][3];
              muxOutConnector[9] = fifoOut[5][3];
              muxOutConnector[10] = fifoOut[6][3];
              muxOutConnector[11] = fifoOut[7][3];
              muxOutConnector[12] = fifoOut[8][3];
              muxOutConnector[13] = fifoOut[9][3];
              muxOutConnector[14] = fifoOut[10][3];
              muxOutConnector[15] = fifoOut[11][3];
              muxOutConnector[16] = fifoOut[12][3];
              muxOutConnector[17] = fifoOut[13][3];
              muxOutConnector[18] = fifoOut[14][3];
              muxOutConnector[19] = fifoOut[15][3];
              muxOutConnector[20] = fifoOut[16][3];
              muxOutConnector[21] = fifoOut[35][0];
              muxOutConnector[22] = fifoOut[36][0];
              muxOutConnector[23] = fifoOut[37][0];
              muxOutConnector[24] = fifoOut[38][0];
              muxOutConnector[25] = fifoOut[39][0];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[17][16];
              muxOutConnector[45] = fifoOut[18][16];
              muxOutConnector[46] = fifoOut[19][16];
              muxOutConnector[47] = fifoOut[20][16];
              muxOutConnector[48] = fifoOut[21][16];
              muxOutConnector[49] = fifoOut[22][16];
              muxOutConnector[50] = fifoOut[23][16];
              muxOutConnector[51] = fifoOut[24][16];
         end
         4: begin
              muxOutConnector[0] = fifoOut[40][1];
              muxOutConnector[1] = fifoOut[41][1];
              muxOutConnector[2] = fifoOut[42][1];
              muxOutConnector[3] = fifoOut[43][1];
              muxOutConnector[4] = fifoOut[44][1];
              muxOutConnector[5] = fifoOut[45][1];
              muxOutConnector[6] = fifoOut[46][1];
              muxOutConnector[7] = fifoOut[47][1];
              muxOutConnector[8] = fifoOut[48][1];
              muxOutConnector[9] = fifoOut[49][1];
              muxOutConnector[10] = fifoOut[50][1];
              muxOutConnector[11] = fifoOut[51][1];
              muxOutConnector[12] = fifoOut[26][0];
              muxOutConnector[13] = fifoOut[27][0];
              muxOutConnector[14] = fifoOut[28][0];
              muxOutConnector[15] = fifoOut[29][0];
              muxOutConnector[16] = fifoOut[30][0];
              muxOutConnector[17] = fifoOut[31][0];
              muxOutConnector[18] = fifoOut[32][0];
              muxOutConnector[19] = fifoOut[33][0];
              muxOutConnector[20] = fifoOut[34][0];
              muxOutConnector[21] = fifoOut[35][0];
              muxOutConnector[22] = fifoOut[36][0];
              muxOutConnector[23] = fifoOut[37][0];
              muxOutConnector[24] = fifoOut[38][0];
              muxOutConnector[25] = fifoOut[39][0];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[17][16];
              muxOutConnector[45] = fifoOut[18][16];
              muxOutConnector[46] = fifoOut[19][16];
              muxOutConnector[47] = fifoOut[20][16];
              muxOutConnector[48] = fifoOut[21][16];
              muxOutConnector[49] = fifoOut[22][16];
              muxOutConnector[50] = fifoOut[23][16];
              muxOutConnector[51] = fifoOut[24][16];
         end
         5: begin
              muxOutConnector[0] = fifoOut[40][1];
              muxOutConnector[1] = fifoOut[41][1];
              muxOutConnector[2] = fifoOut[42][1];
              muxOutConnector[3] = fifoOut[43][1];
              muxOutConnector[4] = fifoOut[44][1];
              muxOutConnector[5] = fifoOut[45][1];
              muxOutConnector[6] = fifoOut[46][1];
              muxOutConnector[7] = fifoOut[47][1];
              muxOutConnector[8] = fifoOut[48][1];
              muxOutConnector[9] = fifoOut[49][1];
              muxOutConnector[10] = fifoOut[50][1];
              muxOutConnector[11] = fifoOut[51][1];
              muxOutConnector[12] = fifoOut[26][0];
              muxOutConnector[13] = fifoOut[27][0];
              muxOutConnector[14] = fifoOut[28][0];
              muxOutConnector[15] = fifoOut[29][0];
              muxOutConnector[16] = fifoOut[30][0];
              muxOutConnector[17] = fifoOut[31][0];
              muxOutConnector[18] = fifoOut[32][0];
              muxOutConnector[19] = fifoOut[33][0];
              muxOutConnector[20] = fifoOut[34][0];
              muxOutConnector[21] = fifoOut[35][0];
              muxOutConnector[22] = fifoOut[36][0];
              muxOutConnector[23] = fifoOut[37][0];
              muxOutConnector[24] = fifoOut[38][0];
              muxOutConnector[25] = fifoOut[39][0];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[17][16];
              muxOutConnector[45] = fifoOut[18][16];
              muxOutConnector[46] = fifoOut[19][16];
              muxOutConnector[47] = fifoOut[20][16];
              muxOutConnector[48] = fifoOut[21][16];
              muxOutConnector[49] = fifoOut[22][16];
              muxOutConnector[50] = fifoOut[23][16];
              muxOutConnector[51] = fifoOut[24][16];
         end
         6: begin
              muxOutConnector[0] = fifoOut[40][1];
              muxOutConnector[1] = fifoOut[41][1];
              muxOutConnector[2] = fifoOut[42][1];
              muxOutConnector[3] = fifoOut[43][1];
              muxOutConnector[4] = fifoOut[44][1];
              muxOutConnector[5] = fifoOut[45][1];
              muxOutConnector[6] = fifoOut[46][1];
              muxOutConnector[7] = fifoOut[47][1];
              muxOutConnector[8] = fifoOut[48][1];
              muxOutConnector[9] = fifoOut[49][1];
              muxOutConnector[10] = fifoOut[50][1];
              muxOutConnector[11] = fifoOut[51][1];
              muxOutConnector[12] = fifoOut[26][0];
              muxOutConnector[13] = fifoOut[27][0];
              muxOutConnector[14] = fifoOut[28][0];
              muxOutConnector[15] = fifoOut[29][0];
              muxOutConnector[16] = fifoOut[30][0];
              muxOutConnector[17] = fifoOut[31][0];
              muxOutConnector[18] = fifoOut[32][0];
              muxOutConnector[19] = fifoOut[33][0];
              muxOutConnector[20] = fifoOut[34][0];
              muxOutConnector[21] = fifoOut[35][0];
              muxOutConnector[22] = fifoOut[36][0];
              muxOutConnector[23] = fifoOut[37][0];
              muxOutConnector[24] = fifoOut[38][0];
              muxOutConnector[25] = fifoOut[39][0];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[17][16];
              muxOutConnector[45] = fifoOut[18][16];
              muxOutConnector[46] = fifoOut[19][16];
              muxOutConnector[47] = fifoOut[20][16];
              muxOutConnector[48] = fifoOut[21][16];
              muxOutConnector[49] = fifoOut[22][16];
              muxOutConnector[50] = fifoOut[23][16];
              muxOutConnector[51] = fifoOut[24][16];
         end
         7: begin
              muxOutConnector[0] = fifoOut[40][1];
              muxOutConnector[1] = fifoOut[41][1];
              muxOutConnector[2] = fifoOut[42][1];
              muxOutConnector[3] = fifoOut[43][1];
              muxOutConnector[4] = fifoOut[44][1];
              muxOutConnector[5] = fifoOut[45][1];
              muxOutConnector[6] = fifoOut[46][1];
              muxOutConnector[7] = fifoOut[47][1];
              muxOutConnector[8] = fifoOut[48][1];
              muxOutConnector[9] = fifoOut[49][1];
              muxOutConnector[10] = fifoOut[50][1];
              muxOutConnector[11] = fifoOut[51][1];
              muxOutConnector[12] = fifoOut[26][0];
              muxOutConnector[13] = fifoOut[27][0];
              muxOutConnector[14] = fifoOut[28][0];
              muxOutConnector[15] = fifoOut[29][0];
              muxOutConnector[16] = fifoOut[30][0];
              muxOutConnector[17] = fifoOut[31][0];
              muxOutConnector[18] = fifoOut[32][0];
              muxOutConnector[19] = fifoOut[33][0];
              muxOutConnector[20] = fifoOut[34][0];
              muxOutConnector[21] = fifoOut[35][0];
              muxOutConnector[22] = fifoOut[36][0];
              muxOutConnector[23] = fifoOut[37][0];
              muxOutConnector[24] = fifoOut[38][0];
              muxOutConnector[25] = fifoOut[39][0];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[17][16];
              muxOutConnector[45] = fifoOut[18][16];
              muxOutConnector[46] = fifoOut[19][16];
              muxOutConnector[47] = fifoOut[20][16];
              muxOutConnector[48] = fifoOut[21][16];
              muxOutConnector[49] = fifoOut[22][16];
              muxOutConnector[50] = fifoOut[23][16];
              muxOutConnector[51] = fifoOut[24][16];
         end
         8: begin
              muxOutConnector[0] = fifoOut[40][1];
              muxOutConnector[1] = fifoOut[41][1];
              muxOutConnector[2] = fifoOut[42][1];
              muxOutConnector[3] = fifoOut[43][1];
              muxOutConnector[4] = fifoOut[44][1];
              muxOutConnector[5] = fifoOut[45][1];
              muxOutConnector[6] = fifoOut[46][1];
              muxOutConnector[7] = fifoOut[47][1];
              muxOutConnector[8] = fifoOut[48][1];
              muxOutConnector[9] = fifoOut[49][1];
              muxOutConnector[10] = fifoOut[50][1];
              muxOutConnector[11] = fifoOut[51][1];
              muxOutConnector[12] = fifoOut[26][0];
              muxOutConnector[13] = fifoOut[27][0];
              muxOutConnector[14] = fifoOut[28][0];
              muxOutConnector[15] = fifoOut[29][0];
              muxOutConnector[16] = fifoOut[30][0];
              muxOutConnector[17] = fifoOut[31][0];
              muxOutConnector[18] = fifoOut[32][0];
              muxOutConnector[19] = fifoOut[33][0];
              muxOutConnector[20] = fifoOut[34][0];
              muxOutConnector[21] = fifoOut[0][5];
              muxOutConnector[22] = fifoOut[1][5];
              muxOutConnector[23] = fifoOut[2][5];
              muxOutConnector[24] = fifoOut[3][5];
              muxOutConnector[25] = fifoOut[4][5];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[17][16];
              muxOutConnector[45] = fifoOut[18][16];
              muxOutConnector[46] = fifoOut[19][16];
              muxOutConnector[47] = fifoOut[20][16];
              muxOutConnector[48] = fifoOut[21][16];
              muxOutConnector[49] = fifoOut[22][16];
              muxOutConnector[50] = fifoOut[23][16];
              muxOutConnector[51] = fifoOut[24][16];
         end
         9: begin
              muxOutConnector[0] = fifoOut[5][6];
              muxOutConnector[1] = fifoOut[6][6];
              muxOutConnector[2] = fifoOut[7][6];
              muxOutConnector[3] = fifoOut[8][6];
              muxOutConnector[4] = fifoOut[9][6];
              muxOutConnector[5] = fifoOut[10][6];
              muxOutConnector[6] = fifoOut[11][6];
              muxOutConnector[7] = fifoOut[12][6];
              muxOutConnector[8] = fifoOut[13][6];
              muxOutConnector[9] = fifoOut[14][6];
              muxOutConnector[10] = fifoOut[15][6];
              muxOutConnector[11] = fifoOut[16][6];
              muxOutConnector[12] = fifoOut[17][6];
              muxOutConnector[13] = fifoOut[18][6];
              muxOutConnector[14] = fifoOut[19][6];
              muxOutConnector[15] = fifoOut[20][6];
              muxOutConnector[16] = fifoOut[21][6];
              muxOutConnector[17] = fifoOut[22][6];
              muxOutConnector[18] = fifoOut[23][6];
              muxOutConnector[19] = fifoOut[24][6];
              muxOutConnector[20] = fifoOut[25][6];
              muxOutConnector[21] = fifoOut[0][5];
              muxOutConnector[22] = fifoOut[1][5];
              muxOutConnector[23] = fifoOut[2][5];
              muxOutConnector[24] = fifoOut[3][5];
              muxOutConnector[25] = fifoOut[4][5];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[17][16];
              muxOutConnector[45] = fifoOut[18][16];
              muxOutConnector[46] = fifoOut[19][16];
              muxOutConnector[47] = fifoOut[20][16];
              muxOutConnector[48] = fifoOut[21][16];
              muxOutConnector[49] = fifoOut[22][16];
              muxOutConnector[50] = fifoOut[23][16];
              muxOutConnector[51] = fifoOut[24][16];
         end
         10: begin
              muxOutConnector[0] = fifoOut[5][6];
              muxOutConnector[1] = fifoOut[6][6];
              muxOutConnector[2] = fifoOut[7][6];
              muxOutConnector[3] = fifoOut[8][6];
              muxOutConnector[4] = fifoOut[9][6];
              muxOutConnector[5] = fifoOut[10][6];
              muxOutConnector[6] = fifoOut[11][6];
              muxOutConnector[7] = fifoOut[12][6];
              muxOutConnector[8] = fifoOut[13][6];
              muxOutConnector[9] = fifoOut[14][6];
              muxOutConnector[10] = fifoOut[15][6];
              muxOutConnector[11] = fifoOut[16][6];
              muxOutConnector[12] = fifoOut[17][6];
              muxOutConnector[13] = fifoOut[18][6];
              muxOutConnector[14] = fifoOut[19][6];
              muxOutConnector[15] = fifoOut[20][6];
              muxOutConnector[16] = fifoOut[21][6];
              muxOutConnector[17] = fifoOut[22][6];
              muxOutConnector[18] = fifoOut[23][6];
              muxOutConnector[19] = fifoOut[24][6];
              muxOutConnector[20] = fifoOut[25][6];
              muxOutConnector[21] = fifoOut[0][5];
              muxOutConnector[22] = fifoOut[1][5];
              muxOutConnector[23] = fifoOut[2][5];
              muxOutConnector[24] = fifoOut[3][5];
              muxOutConnector[25] = fifoOut[4][5];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[17][16];
              muxOutConnector[45] = fifoOut[18][16];
              muxOutConnector[46] = fifoOut[19][16];
              muxOutConnector[47] = fifoOut[20][16];
              muxOutConnector[48] = fifoOut[21][16];
              muxOutConnector[49] = fifoOut[22][16];
              muxOutConnector[50] = fifoOut[23][16];
              muxOutConnector[51] = fifoOut[24][16];
         end
         11: begin
              muxOutConnector[0] = fifoOut[5][6];
              muxOutConnector[1] = fifoOut[6][6];
              muxOutConnector[2] = fifoOut[7][6];
              muxOutConnector[3] = fifoOut[8][6];
              muxOutConnector[4] = fifoOut[9][6];
              muxOutConnector[5] = fifoOut[10][6];
              muxOutConnector[6] = fifoOut[11][6];
              muxOutConnector[7] = fifoOut[12][6];
              muxOutConnector[8] = fifoOut[13][6];
              muxOutConnector[9] = fifoOut[14][6];
              muxOutConnector[10] = fifoOut[15][6];
              muxOutConnector[11] = fifoOut[16][6];
              muxOutConnector[12] = fifoOut[17][6];
              muxOutConnector[13] = fifoOut[18][6];
              muxOutConnector[14] = fifoOut[19][6];
              muxOutConnector[15] = fifoOut[20][6];
              muxOutConnector[16] = fifoOut[21][6];
              muxOutConnector[17] = fifoOut[22][6];
              muxOutConnector[18] = fifoOut[23][6];
              muxOutConnector[19] = fifoOut[24][6];
              muxOutConnector[20] = fifoOut[25][6];
              muxOutConnector[21] = fifoOut[0][5];
              muxOutConnector[22] = fifoOut[1][5];
              muxOutConnector[23] = fifoOut[2][5];
              muxOutConnector[24] = fifoOut[3][5];
              muxOutConnector[25] = fifoOut[4][5];
              muxOutConnector[26] = fifoOut[34][11];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[17][16];
              muxOutConnector[45] = fifoOut[18][16];
              muxOutConnector[46] = fifoOut[19][16];
              muxOutConnector[47] = fifoOut[20][16];
              muxOutConnector[48] = fifoOut[21][16];
              muxOutConnector[49] = fifoOut[22][16];
              muxOutConnector[50] = fifoOut[23][16];
              muxOutConnector[51] = fifoOut[24][16];
         end
         12: begin
              muxOutConnector[0] = fifoOut[5][6];
              muxOutConnector[1] = fifoOut[6][6];
              muxOutConnector[2] = fifoOut[7][6];
              muxOutConnector[3] = fifoOut[8][6];
              muxOutConnector[4] = fifoOut[9][6];
              muxOutConnector[5] = fifoOut[10][6];
              muxOutConnector[6] = fifoOut[11][6];
              muxOutConnector[7] = fifoOut[12][6];
              muxOutConnector[8] = fifoOut[13][6];
              muxOutConnector[9] = fifoOut[14][6];
              muxOutConnector[10] = fifoOut[15][6];
              muxOutConnector[11] = fifoOut[16][6];
              muxOutConnector[12] = fifoOut[17][6];
              muxOutConnector[13] = fifoOut[18][6];
              muxOutConnector[14] = fifoOut[19][6];
              muxOutConnector[15] = fifoOut[20][6];
              muxOutConnector[16] = fifoOut[21][6];
              muxOutConnector[17] = fifoOut[22][6];
              muxOutConnector[18] = fifoOut[23][6];
              muxOutConnector[19] = fifoOut[24][6];
              muxOutConnector[20] = fifoOut[25][6];
              muxOutConnector[21] = fifoOut[0][5];
              muxOutConnector[22] = fifoOut[1][5];
              muxOutConnector[23] = fifoOut[2][5];
              muxOutConnector[24] = fifoOut[3][5];
              muxOutConnector[25] = fifoOut[4][5];
              muxOutConnector[26] = fifoOut[25][0];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[17][16];
              muxOutConnector[45] = fifoOut[18][16];
              muxOutConnector[46] = fifoOut[19][16];
              muxOutConnector[47] = fifoOut[20][16];
              muxOutConnector[48] = fifoOut[21][16];
              muxOutConnector[49] = fifoOut[22][16];
              muxOutConnector[50] = fifoOut[23][16];
              muxOutConnector[51] = fifoOut[24][16];
         end
         13: begin
              muxOutConnector[0] = fifoOut[5][6];
              muxOutConnector[1] = fifoOut[6][6];
              muxOutConnector[2] = fifoOut[7][6];
              muxOutConnector[3] = fifoOut[8][6];
              muxOutConnector[4] = fifoOut[9][6];
              muxOutConnector[5] = fifoOut[10][6];
              muxOutConnector[6] = fifoOut[11][6];
              muxOutConnector[7] = fifoOut[12][6];
              muxOutConnector[8] = fifoOut[13][6];
              muxOutConnector[9] = fifoOut[14][6];
              muxOutConnector[10] = fifoOut[15][6];
              muxOutConnector[11] = fifoOut[16][6];
              muxOutConnector[12] = fifoOut[17][6];
              muxOutConnector[13] = fifoOut[18][6];
              muxOutConnector[14] = fifoOut[19][6];
              muxOutConnector[15] = fifoOut[20][6];
              muxOutConnector[16] = fifoOut[21][6];
              muxOutConnector[17] = fifoOut[22][6];
              muxOutConnector[18] = fifoOut[23][6];
              muxOutConnector[19] = fifoOut[24][6];
              muxOutConnector[20] = fifoOut[25][6];
              muxOutConnector[21] = fifoOut[0][5];
              muxOutConnector[22] = fifoOut[1][5];
              muxOutConnector[23] = fifoOut[2][5];
              muxOutConnector[24] = fifoOut[3][5];
              muxOutConnector[25] = fifoOut[4][5];
              muxOutConnector[26] = fifoOut[25][0];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[17][16];
              muxOutConnector[45] = fifoOut[18][16];
              muxOutConnector[46] = fifoOut[19][16];
              muxOutConnector[47] = fifoOut[20][16];
              muxOutConnector[48] = fifoOut[21][16];
              muxOutConnector[49] = fifoOut[22][16];
              muxOutConnector[50] = fifoOut[23][16];
              muxOutConnector[51] = fifoOut[24][16];
         end
         14: begin
              muxOutConnector[0] = fifoOut[5][6];
              muxOutConnector[1] = fifoOut[6][6];
              muxOutConnector[2] = fifoOut[7][6];
              muxOutConnector[3] = fifoOut[8][6];
              muxOutConnector[4] = fifoOut[9][6];
              muxOutConnector[5] = fifoOut[10][6];
              muxOutConnector[6] = fifoOut[11][6];
              muxOutConnector[7] = fifoOut[12][6];
              muxOutConnector[8] = fifoOut[13][6];
              muxOutConnector[9] = fifoOut[14][6];
              muxOutConnector[10] = fifoOut[15][6];
              muxOutConnector[11] = fifoOut[16][6];
              muxOutConnector[12] = fifoOut[17][6];
              muxOutConnector[13] = fifoOut[18][6];
              muxOutConnector[14] = fifoOut[19][6];
              muxOutConnector[15] = fifoOut[20][6];
              muxOutConnector[16] = fifoOut[21][6];
              muxOutConnector[17] = fifoOut[22][6];
              muxOutConnector[18] = fifoOut[23][6];
              muxOutConnector[19] = fifoOut[24][6];
              muxOutConnector[20] = fifoOut[25][6];
              muxOutConnector[21] = fifoOut[0][5];
              muxOutConnector[22] = fifoOut[1][5];
              muxOutConnector[23] = fifoOut[2][5];
              muxOutConnector[24] = fifoOut[3][5];
              muxOutConnector[25] = fifoOut[4][5];
              muxOutConnector[26] = fifoOut[25][0];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[17][16];
              muxOutConnector[45] = fifoOut[18][16];
              muxOutConnector[46] = fifoOut[19][16];
              muxOutConnector[47] = fifoOut[20][16];
              muxOutConnector[48] = fifoOut[21][16];
              muxOutConnector[49] = fifoOut[22][16];
              muxOutConnector[50] = fifoOut[23][16];
              muxOutConnector[51] = fifoOut[24][16];
         end
         15: begin
              muxOutConnector[0] = fifoOut[5][6];
              muxOutConnector[1] = fifoOut[6][6];
              muxOutConnector[2] = fifoOut[7][6];
              muxOutConnector[3] = fifoOut[8][6];
              muxOutConnector[4] = fifoOut[9][6];
              muxOutConnector[5] = fifoOut[10][6];
              muxOutConnector[6] = fifoOut[11][6];
              muxOutConnector[7] = fifoOut[12][6];
              muxOutConnector[8] = fifoOut[13][6];
              muxOutConnector[9] = fifoOut[14][6];
              muxOutConnector[10] = fifoOut[15][6];
              muxOutConnector[11] = fifoOut[16][6];
              muxOutConnector[12] = fifoOut[17][6];
              muxOutConnector[13] = fifoOut[18][6];
              muxOutConnector[14] = fifoOut[19][6];
              muxOutConnector[15] = fifoOut[20][6];
              muxOutConnector[16] = fifoOut[21][6];
              muxOutConnector[17] = fifoOut[22][6];
              muxOutConnector[18] = fifoOut[23][6];
              muxOutConnector[19] = fifoOut[24][6];
              muxOutConnector[20] = fifoOut[25][6];
              muxOutConnector[21] = fifoOut[0][5];
              muxOutConnector[22] = fifoOut[1][5];
              muxOutConnector[23] = fifoOut[2][5];
              muxOutConnector[24] = fifoOut[3][5];
              muxOutConnector[25] = fifoOut[4][5];
              muxOutConnector[26] = fifoOut[25][0];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[17][16];
              muxOutConnector[45] = fifoOut[18][16];
              muxOutConnector[46] = fifoOut[19][16];
              muxOutConnector[47] = fifoOut[20][16];
              muxOutConnector[48] = fifoOut[21][16];
              muxOutConnector[49] = fifoOut[22][16];
              muxOutConnector[50] = fifoOut[23][16];
              muxOutConnector[51] = fifoOut[24][16];
         end
         16: begin
              muxOutConnector[0] = fifoOut[5][6];
              muxOutConnector[1] = fifoOut[6][6];
              muxOutConnector[2] = fifoOut[7][6];
              muxOutConnector[3] = fifoOut[8][6];
              muxOutConnector[4] = fifoOut[9][6];
              muxOutConnector[5] = fifoOut[10][6];
              muxOutConnector[6] = fifoOut[11][6];
              muxOutConnector[7] = fifoOut[12][6];
              muxOutConnector[8] = fifoOut[13][6];
              muxOutConnector[9] = fifoOut[14][6];
              muxOutConnector[10] = fifoOut[15][6];
              muxOutConnector[11] = fifoOut[16][6];
              muxOutConnector[12] = fifoOut[17][6];
              muxOutConnector[13] = fifoOut[18][6];
              muxOutConnector[14] = fifoOut[19][6];
              muxOutConnector[15] = fifoOut[20][6];
              muxOutConnector[16] = fifoOut[21][6];
              muxOutConnector[17] = fifoOut[22][6];
              muxOutConnector[18] = fifoOut[23][6];
              muxOutConnector[19] = fifoOut[24][6];
              muxOutConnector[20] = fifoOut[25][6];
              muxOutConnector[21] = fifoOut[0][5];
              muxOutConnector[22] = fifoOut[1][5];
              muxOutConnector[23] = fifoOut[2][5];
              muxOutConnector[24] = fifoOut[3][5];
              muxOutConnector[25] = fifoOut[4][5];
              muxOutConnector[26] = fifoOut[25][0];
              muxOutConnector[27] = fifoOut[0][16];
              muxOutConnector[28] = fifoOut[1][16];
              muxOutConnector[29] = fifoOut[2][16];
              muxOutConnector[30] = fifoOut[3][16];
              muxOutConnector[31] = fifoOut[4][16];
              muxOutConnector[32] = fifoOut[5][16];
              muxOutConnector[33] = fifoOut[6][16];
              muxOutConnector[34] = fifoOut[7][16];
              muxOutConnector[35] = fifoOut[8][16];
              muxOutConnector[36] = fifoOut[9][16];
              muxOutConnector[37] = fifoOut[10][16];
              muxOutConnector[38] = fifoOut[11][16];
              muxOutConnector[39] = fifoOut[12][16];
              muxOutConnector[40] = fifoOut[13][16];
              muxOutConnector[41] = fifoOut[14][16];
              muxOutConnector[42] = fifoOut[15][16];
              muxOutConnector[43] = fifoOut[16][16];
              muxOutConnector[44] = fifoOut[35][13];
              muxOutConnector[45] = fifoOut[36][13];
              muxOutConnector[46] = fifoOut[37][13];
              muxOutConnector[47] = fifoOut[38][13];
              muxOutConnector[48] = fifoOut[39][13];
              muxOutConnector[49] = fifoOut[40][13];
              muxOutConnector[50] = fifoOut[41][13];
              muxOutConnector[51] = fifoOut[42][13];
         end
         17: begin
              muxOutConnector[0] = fifoOut[5][6];
              muxOutConnector[1] = fifoOut[6][6];
              muxOutConnector[2] = fifoOut[7][6];
              muxOutConnector[3] = fifoOut[8][6];
              muxOutConnector[4] = fifoOut[9][6];
              muxOutConnector[5] = fifoOut[10][6];
              muxOutConnector[6] = fifoOut[11][6];
              muxOutConnector[7] = fifoOut[12][6];
              muxOutConnector[8] = fifoOut[13][6];
              muxOutConnector[9] = fifoOut[14][6];
              muxOutConnector[10] = fifoOut[15][6];
              muxOutConnector[11] = fifoOut[16][6];
              muxOutConnector[12] = fifoOut[17][6];
              muxOutConnector[13] = fifoOut[18][6];
              muxOutConnector[14] = fifoOut[19][6];
              muxOutConnector[15] = fifoOut[20][6];
              muxOutConnector[16] = fifoOut[21][6];
              muxOutConnector[17] = fifoOut[22][6];
              muxOutConnector[18] = fifoOut[23][6];
              muxOutConnector[19] = fifoOut[24][6];
              muxOutConnector[20] = fifoOut[25][6];
              muxOutConnector[21] = fifoOut[0][5];
              muxOutConnector[22] = fifoOut[1][5];
              muxOutConnector[23] = fifoOut[2][5];
              muxOutConnector[24] = fifoOut[3][5];
              muxOutConnector[25] = fifoOut[4][5];
              muxOutConnector[26] = fifoOut[43][14];
              muxOutConnector[27] = fifoOut[44][14];
              muxOutConnector[28] = fifoOut[45][14];
              muxOutConnector[29] = fifoOut[46][14];
              muxOutConnector[30] = fifoOut[47][14];
              muxOutConnector[31] = fifoOut[48][14];
              muxOutConnector[32] = fifoOut[49][14];
              muxOutConnector[33] = fifoOut[50][14];
              muxOutConnector[34] = fifoOut[51][14];
              muxOutConnector[35] = fifoOut[26][13];
              muxOutConnector[36] = fifoOut[27][13];
              muxOutConnector[37] = fifoOut[28][13];
              muxOutConnector[38] = fifoOut[29][13];
              muxOutConnector[39] = fifoOut[30][13];
              muxOutConnector[40] = fifoOut[31][13];
              muxOutConnector[41] = fifoOut[32][13];
              muxOutConnector[42] = fifoOut[33][13];
              muxOutConnector[43] = fifoOut[34][13];
              muxOutConnector[44] = fifoOut[35][13];
              muxOutConnector[45] = fifoOut[36][13];
              muxOutConnector[46] = fifoOut[37][13];
              muxOutConnector[47] = fifoOut[38][13];
              muxOutConnector[48] = fifoOut[39][13];
              muxOutConnector[49] = fifoOut[40][13];
              muxOutConnector[50] = fifoOut[41][13];
              muxOutConnector[51] = fifoOut[42][13];
         end
         18: begin
              muxOutConnector[0] = fifoOut[5][6];
              muxOutConnector[1] = fifoOut[6][6];
              muxOutConnector[2] = fifoOut[7][6];
              muxOutConnector[3] = fifoOut[8][6];
              muxOutConnector[4] = fifoOut[9][6];
              muxOutConnector[5] = fifoOut[10][6];
              muxOutConnector[6] = fifoOut[11][6];
              muxOutConnector[7] = fifoOut[12][6];
              muxOutConnector[8] = fifoOut[13][6];
              muxOutConnector[9] = fifoOut[14][6];
              muxOutConnector[10] = fifoOut[15][6];
              muxOutConnector[11] = fifoOut[16][6];
              muxOutConnector[12] = fifoOut[17][6];
              muxOutConnector[13] = fifoOut[18][6];
              muxOutConnector[14] = fifoOut[19][6];
              muxOutConnector[15] = fifoOut[20][6];
              muxOutConnector[16] = fifoOut[21][6];
              muxOutConnector[17] = fifoOut[22][6];
              muxOutConnector[18] = fifoOut[23][6];
              muxOutConnector[19] = fifoOut[24][6];
              muxOutConnector[20] = fifoOut[25][6];
              muxOutConnector[21] = fifoOut[0][5];
              muxOutConnector[22] = fifoOut[1][5];
              muxOutConnector[23] = fifoOut[2][5];
              muxOutConnector[24] = fifoOut[3][5];
              muxOutConnector[25] = fifoOut[4][5];
              muxOutConnector[26] = fifoOut[43][14];
              muxOutConnector[27] = fifoOut[44][14];
              muxOutConnector[28] = fifoOut[45][14];
              muxOutConnector[29] = fifoOut[46][14];
              muxOutConnector[30] = fifoOut[47][14];
              muxOutConnector[31] = fifoOut[48][14];
              muxOutConnector[32] = fifoOut[49][14];
              muxOutConnector[33] = fifoOut[50][14];
              muxOutConnector[34] = fifoOut[51][14];
              muxOutConnector[35] = fifoOut[26][13];
              muxOutConnector[36] = fifoOut[27][13];
              muxOutConnector[37] = fifoOut[28][13];
              muxOutConnector[38] = fifoOut[29][13];
              muxOutConnector[39] = fifoOut[30][13];
              muxOutConnector[40] = fifoOut[31][13];
              muxOutConnector[41] = fifoOut[32][13];
              muxOutConnector[42] = fifoOut[33][13];
              muxOutConnector[43] = fifoOut[34][13];
              muxOutConnector[44] = fifoOut[35][13];
              muxOutConnector[45] = fifoOut[36][13];
              muxOutConnector[46] = fifoOut[37][13];
              muxOutConnector[47] = fifoOut[38][13];
              muxOutConnector[48] = fifoOut[39][13];
              muxOutConnector[49] = fifoOut[40][13];
              muxOutConnector[50] = fifoOut[41][13];
              muxOutConnector[51] = fifoOut[42][13];
         end
         19: begin
              muxOutConnector[0] = fifoOut[5][6];
              muxOutConnector[1] = fifoOut[6][6];
              muxOutConnector[2] = fifoOut[7][6];
              muxOutConnector[3] = fifoOut[8][6];
              muxOutConnector[4] = fifoOut[9][6];
              muxOutConnector[5] = fifoOut[10][6];
              muxOutConnector[6] = fifoOut[11][6];
              muxOutConnector[7] = fifoOut[12][6];
              muxOutConnector[8] = fifoOut[13][6];
              muxOutConnector[9] = fifoOut[14][6];
              muxOutConnector[10] = fifoOut[15][6];
              muxOutConnector[11] = fifoOut[16][6];
              muxOutConnector[12] = fifoOut[17][6];
              muxOutConnector[13] = fifoOut[18][6];
              muxOutConnector[14] = fifoOut[19][6];
              muxOutConnector[15] = fifoOut[20][6];
              muxOutConnector[16] = fifoOut[21][6];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[43][14];
              muxOutConnector[27] = fifoOut[44][14];
              muxOutConnector[28] = fifoOut[45][14];
              muxOutConnector[29] = fifoOut[46][14];
              muxOutConnector[30] = fifoOut[47][14];
              muxOutConnector[31] = fifoOut[48][14];
              muxOutConnector[32] = fifoOut[49][14];
              muxOutConnector[33] = fifoOut[50][14];
              muxOutConnector[34] = fifoOut[51][14];
              muxOutConnector[35] = fifoOut[26][13];
              muxOutConnector[36] = fifoOut[27][13];
              muxOutConnector[37] = fifoOut[28][13];
              muxOutConnector[38] = fifoOut[29][13];
              muxOutConnector[39] = fifoOut[30][13];
              muxOutConnector[40] = fifoOut[31][13];
              muxOutConnector[41] = fifoOut[32][13];
              muxOutConnector[42] = fifoOut[33][13];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
         end
         default: begin
               for(i=0;i<muxOutSymbols;i=i+1)begin
                muxOutConnector[i] = 0;
              end
         end
//hgjhgbuiguigbigbgbgbui
         endcase
    end
       1: begin // iteration_0_indicator = 0
    case(rd_address_case)
      0: begin
           muxOutConnector[0] = maxVal;
           muxOutConnector[1] = maxVal;
           muxOutConnector[2] = maxVal;
           muxOutConnector[3] = maxVal;
           muxOutConnector[4] = maxVal;
           muxOutConnector[5] = maxVal;
           muxOutConnector[6] = maxVal;
           muxOutConnector[7] = maxVal;
           muxOutConnector[8] = maxVal;
           muxOutConnector[9] = maxVal;
           muxOutConnector[10] = maxVal;
           muxOutConnector[11] = maxVal;
           muxOutConnector[12] = maxVal;
           muxOutConnector[13] = maxVal;
           muxOutConnector[14] = maxVal;
           muxOutConnector[15] = maxVal;
           muxOutConnector[16] = maxVal;
           muxOutConnector[17] = maxVal;
           muxOutConnector[18] = fifoOut[0][15];
           muxOutConnector[19] = fifoOut[1][15];
           muxOutConnector[20] = fifoOut[2][15];
           muxOutConnector[21] = fifoOut[3][15];
           muxOutConnector[22] = fifoOut[4][15];
           muxOutConnector[23] = fifoOut[5][15];
           muxOutConnector[24] = fifoOut[6][15];
           muxOutConnector[25] = fifoOut[7][15];
           muxOutConnector[26] = fifoOut[30][11];
           muxOutConnector[27] = fifoOut[31][11];
           muxOutConnector[28] = fifoOut[0][10];
           muxOutConnector[29] = fifoOut[1][10];
           muxOutConnector[30] = fifoOut[2][10];
           muxOutConnector[31] = fifoOut[3][10];
           muxOutConnector[32] = fifoOut[4][10];
           muxOutConnector[33] = fifoOut[5][10];
           muxOutConnector[34] = fifoOut[6][10];
           muxOutConnector[35] = fifoOut[7][10];
           muxOutConnector[36] = fifoOut[8][10];
           muxOutConnector[37] = fifoOut[9][10];
           muxOutConnector[38] = fifoOut[10][10];
           muxOutConnector[39] = fifoOut[11][10];
           muxOutConnector[40] = fifoOut[12][10];
           muxOutConnector[41] = fifoOut[13][10];
           muxOutConnector[42] = fifoOut[14][10];
           muxOutConnector[43] = fifoOut[15][10];
           muxOutConnector[44] = fifoOut[16][10];
           muxOutConnector[45] = fifoOut[17][10];
           muxOutConnector[46] = fifoOut[18][10];
           muxOutConnector[47] = fifoOut[19][10];
           muxOutConnector[48] = fifoOut[20][10];
           muxOutConnector[49] = fifoOut[21][10];
           muxOutConnector[50] = fifoOut[22][10];
           muxOutConnector[51] = fifoOut[23][10];
      end
      1: begin
           muxOutConnector[0] = fifoOut[8][16];
           muxOutConnector[1] = fifoOut[9][16];
           muxOutConnector[2] = fifoOut[10][16];
           muxOutConnector[3] = fifoOut[11][16];
           muxOutConnector[4] = fifoOut[12][16];
           muxOutConnector[5] = fifoOut[13][16];
           muxOutConnector[6] = fifoOut[14][16];
           muxOutConnector[7] = fifoOut[15][16];
           muxOutConnector[8] = fifoOut[16][16];
           muxOutConnector[9] = fifoOut[17][16];
           muxOutConnector[10] = fifoOut[18][16];
           muxOutConnector[11] = fifoOut[19][16];
           muxOutConnector[12] = fifoOut[20][16];
           muxOutConnector[13] = fifoOut[21][16];
           muxOutConnector[14] = fifoOut[22][16];
           muxOutConnector[15] = fifoOut[23][16];
           muxOutConnector[16] = fifoOut[24][16];
           muxOutConnector[17] = fifoOut[25][16];
           muxOutConnector[18] = fifoOut[26][16];
           muxOutConnector[19] = fifoOut[27][16];
           muxOutConnector[20] = fifoOut[28][16];
           muxOutConnector[21] = fifoOut[29][16];
           muxOutConnector[22] = fifoOut[30][16];
           muxOutConnector[23] = fifoOut[31][16];
           muxOutConnector[24] = fifoOut[0][15];
           muxOutConnector[25] = fifoOut[1][15];
           muxOutConnector[26] = fifoOut[24][11];
           muxOutConnector[27] = fifoOut[25][11];
           muxOutConnector[28] = fifoOut[26][11];
           muxOutConnector[29] = fifoOut[27][11];
           muxOutConnector[30] = fifoOut[28][11];
           muxOutConnector[31] = fifoOut[29][11];
           muxOutConnector[32] = fifoOut[30][11];
           muxOutConnector[33] = fifoOut[31][11];
           muxOutConnector[34] = fifoOut[0][10];
           muxOutConnector[35] = fifoOut[1][10];
           muxOutConnector[36] = fifoOut[2][10];
           muxOutConnector[37] = fifoOut[3][10];
           muxOutConnector[38] = fifoOut[4][10];
           muxOutConnector[39] = fifoOut[5][10];
           muxOutConnector[40] = fifoOut[6][10];
           muxOutConnector[41] = fifoOut[7][10];
           muxOutConnector[42] = fifoOut[8][10];
           muxOutConnector[43] = fifoOut[9][10];
           muxOutConnector[44] = fifoOut[10][10];
           muxOutConnector[45] = fifoOut[11][10];
           muxOutConnector[46] = fifoOut[12][10];
           muxOutConnector[47] = fifoOut[13][10];
           muxOutConnector[48] = fifoOut[14][10];
           muxOutConnector[49] = fifoOut[15][10];
           muxOutConnector[50] = fifoOut[16][10];
           muxOutConnector[51] = fifoOut[17][10];
      end
      2: begin
           muxOutConnector[0] = fifoOut[2][16];
           muxOutConnector[1] = fifoOut[3][16];
           muxOutConnector[2] = fifoOut[4][16];
           muxOutConnector[3] = fifoOut[5][16];
           muxOutConnector[4] = fifoOut[6][16];
           muxOutConnector[5] = fifoOut[7][16];
           muxOutConnector[6] = fifoOut[8][16];
           muxOutConnector[7] = fifoOut[9][16];
           muxOutConnector[8] = fifoOut[10][16];
           muxOutConnector[9] = fifoOut[11][16];
           muxOutConnector[10] = fifoOut[12][16];
           muxOutConnector[11] = fifoOut[13][16];
           muxOutConnector[12] = fifoOut[14][16];
           muxOutConnector[13] = fifoOut[15][16];
           muxOutConnector[14] = fifoOut[16][16];
           muxOutConnector[15] = fifoOut[17][16];
           muxOutConnector[16] = fifoOut[18][16];
           muxOutConnector[17] = fifoOut[19][16];
           muxOutConnector[18] = fifoOut[20][16];
           muxOutConnector[19] = fifoOut[21][16];
           muxOutConnector[20] = fifoOut[22][16];
           muxOutConnector[21] = fifoOut[23][16];
           muxOutConnector[22] = fifoOut[24][16];
           muxOutConnector[23] = fifoOut[25][16];
           muxOutConnector[24] = fifoOut[26][16];
           muxOutConnector[25] = fifoOut[27][16];
           muxOutConnector[26] = fifoOut[18][11];
           muxOutConnector[27] = fifoOut[19][11];
           muxOutConnector[28] = fifoOut[20][11];
           muxOutConnector[29] = fifoOut[21][11];
           muxOutConnector[30] = fifoOut[22][11];
           muxOutConnector[31] = fifoOut[23][11];
           muxOutConnector[32] = fifoOut[24][11];
           muxOutConnector[33] = fifoOut[25][11];
           muxOutConnector[34] = fifoOut[26][11];
           muxOutConnector[35] = fifoOut[27][11];
           muxOutConnector[36] = fifoOut[28][11];
           muxOutConnector[37] = fifoOut[29][11];
           muxOutConnector[38] = fifoOut[30][11];
           muxOutConnector[39] = fifoOut[31][11];
           muxOutConnector[40] = fifoOut[0][10];
           muxOutConnector[41] = fifoOut[1][10];
           muxOutConnector[42] = fifoOut[2][10];
           muxOutConnector[43] = fifoOut[3][10];
           muxOutConnector[44] = fifoOut[4][10];
           muxOutConnector[45] = fifoOut[5][10];
           muxOutConnector[46] = fifoOut[6][10];
           muxOutConnector[47] = fifoOut[7][10];
           muxOutConnector[48] = fifoOut[8][10];
           muxOutConnector[49] = fifoOut[9][10];
           muxOutConnector[50] = fifoOut[10][10];
           muxOutConnector[51] = fifoOut[11][10];
      end
      3: begin
           muxOutConnector[0] = fifoOut[28][0];
           muxOutConnector[1] = fifoOut[29][0];
           muxOutConnector[2] = fifoOut[30][0];
           muxOutConnector[3] = fifoOut[31][0];
           muxOutConnector[4] = fifoOut[0][16];
           muxOutConnector[5] = fifoOut[1][16];
           muxOutConnector[6] = fifoOut[2][16];
           muxOutConnector[7] = fifoOut[3][16];
           muxOutConnector[8] = fifoOut[4][16];
           muxOutConnector[9] = fifoOut[5][16];
           muxOutConnector[10] = fifoOut[6][16];
           muxOutConnector[11] = fifoOut[7][16];
           muxOutConnector[12] = fifoOut[8][16];
           muxOutConnector[13] = fifoOut[9][16];
           muxOutConnector[14] = fifoOut[10][16];
           muxOutConnector[15] = fifoOut[11][16];
           muxOutConnector[16] = fifoOut[12][16];
           muxOutConnector[17] = fifoOut[13][16];
           muxOutConnector[18] = fifoOut[14][16];
           muxOutConnector[19] = fifoOut[15][16];
           muxOutConnector[20] = fifoOut[16][16];
           muxOutConnector[21] = fifoOut[17][16];
           muxOutConnector[22] = fifoOut[18][16];
           muxOutConnector[23] = fifoOut[19][16];
           muxOutConnector[24] = fifoOut[20][16];
           muxOutConnector[25] = fifoOut[21][16];
           muxOutConnector[26] = fifoOut[12][11];
           muxOutConnector[27] = fifoOut[13][11];
           muxOutConnector[28] = fifoOut[14][11];
           muxOutConnector[29] = fifoOut[15][11];
           muxOutConnector[30] = fifoOut[16][11];
           muxOutConnector[31] = fifoOut[17][11];
           muxOutConnector[32] = fifoOut[18][11];
           muxOutConnector[33] = fifoOut[19][11];
           muxOutConnector[34] = fifoOut[20][11];
           muxOutConnector[35] = fifoOut[21][11];
           muxOutConnector[36] = fifoOut[22][11];
           muxOutConnector[37] = fifoOut[23][11];
           muxOutConnector[38] = fifoOut[24][11];
           muxOutConnector[39] = fifoOut[25][11];
           muxOutConnector[40] = fifoOut[26][11];
           muxOutConnector[41] = fifoOut[27][11];
           muxOutConnector[42] = fifoOut[28][11];
           muxOutConnector[43] = fifoOut[29][11];
           muxOutConnector[44] = fifoOut[30][11];
           muxOutConnector[45] = fifoOut[31][11];
           muxOutConnector[46] = fifoOut[0][10];
           muxOutConnector[47] = fifoOut[1][10];
           muxOutConnector[48] = fifoOut[2][10];
           muxOutConnector[49] = fifoOut[3][10];
           muxOutConnector[50] = fifoOut[4][10];
           muxOutConnector[51] = fifoOut[5][10];
      end
      4: begin
           muxOutConnector[0] = fifoOut[22][0];
           muxOutConnector[1] = fifoOut[23][0];
           muxOutConnector[2] = fifoOut[24][0];
           muxOutConnector[3] = fifoOut[25][0];
           muxOutConnector[4] = fifoOut[26][0];
           muxOutConnector[5] = fifoOut[27][0];
           muxOutConnector[6] = fifoOut[28][0];
           muxOutConnector[7] = fifoOut[29][0];
           muxOutConnector[8] = fifoOut[30][0];
           muxOutConnector[9] = fifoOut[31][0];
           muxOutConnector[10] = fifoOut[0][16];
           muxOutConnector[11] = fifoOut[1][16];
           muxOutConnector[12] = fifoOut[2][16];
           muxOutConnector[13] = fifoOut[3][16];
           muxOutConnector[14] = fifoOut[4][16];
           muxOutConnector[15] = fifoOut[5][16];
           muxOutConnector[16] = fifoOut[6][16];
           muxOutConnector[17] = fifoOut[7][16];
           muxOutConnector[18] = fifoOut[8][16];
           muxOutConnector[19] = fifoOut[9][16];
           muxOutConnector[20] = fifoOut[10][16];
           muxOutConnector[21] = fifoOut[11][16];
           muxOutConnector[22] = fifoOut[12][16];
           muxOutConnector[23] = fifoOut[13][16];
           muxOutConnector[24] = fifoOut[14][16];
           muxOutConnector[25] = fifoOut[15][16];
           muxOutConnector[26] = fifoOut[6][11];
           muxOutConnector[27] = fifoOut[7][11];
           muxOutConnector[28] = fifoOut[8][11];
           muxOutConnector[29] = fifoOut[9][11];
           muxOutConnector[30] = fifoOut[10][11];
           muxOutConnector[31] = fifoOut[11][11];
           muxOutConnector[32] = fifoOut[12][11];
           muxOutConnector[33] = fifoOut[13][11];
           muxOutConnector[34] = fifoOut[14][11];
           muxOutConnector[35] = fifoOut[15][11];
           muxOutConnector[36] = fifoOut[16][11];
           muxOutConnector[37] = fifoOut[17][11];
           muxOutConnector[38] = fifoOut[18][11];
           muxOutConnector[39] = fifoOut[19][11];
           muxOutConnector[40] = fifoOut[20][11];
           muxOutConnector[41] = fifoOut[21][11];
           muxOutConnector[42] = fifoOut[22][11];
           muxOutConnector[43] = fifoOut[23][11];
           muxOutConnector[44] = fifoOut[24][11];
           muxOutConnector[45] = fifoOut[25][11];
           muxOutConnector[46] = fifoOut[26][11];
           muxOutConnector[47] = fifoOut[27][11];
           muxOutConnector[48] = fifoOut[28][11];
           muxOutConnector[49] = fifoOut[29][11];
           muxOutConnector[50] = fifoOut[30][11];
           muxOutConnector[51] = fifoOut[31][11];
      end
      5: begin
           muxOutConnector[0] = fifoOut[16][0];
           muxOutConnector[1] = fifoOut[17][0];
           muxOutConnector[2] = fifoOut[18][0];
           muxOutConnector[3] = fifoOut[19][0];
           muxOutConnector[4] = fifoOut[20][0];
           muxOutConnector[5] = fifoOut[21][0];
           muxOutConnector[6] = fifoOut[22][0];
           muxOutConnector[7] = fifoOut[23][0];
           muxOutConnector[8] = fifoOut[24][0];
           muxOutConnector[9] = fifoOut[25][0];
           muxOutConnector[10] = fifoOut[26][0];
           muxOutConnector[11] = fifoOut[27][0];
           muxOutConnector[12] = fifoOut[28][0];
           muxOutConnector[13] = fifoOut[29][0];
           muxOutConnector[14] = fifoOut[30][0];
           muxOutConnector[15] = fifoOut[31][0];
           muxOutConnector[16] = fifoOut[0][16];
           muxOutConnector[17] = fifoOut[1][16];
           muxOutConnector[18] = fifoOut[2][16];
           muxOutConnector[19] = fifoOut[3][16];
           muxOutConnector[20] = fifoOut[4][16];
           muxOutConnector[21] = fifoOut[5][16];
           muxOutConnector[22] = fifoOut[6][16];
           muxOutConnector[23] = fifoOut[7][16];
           muxOutConnector[24] = fifoOut[8][16];
           muxOutConnector[25] = fifoOut[9][16];
           muxOutConnector[26] = fifoOut[0][11];
           muxOutConnector[27] = fifoOut[1][11];
           muxOutConnector[28] = fifoOut[2][11];
           muxOutConnector[29] = fifoOut[3][11];
           muxOutConnector[30] = fifoOut[4][11];
           muxOutConnector[31] = fifoOut[5][11];
           muxOutConnector[32] = fifoOut[6][11];
           muxOutConnector[33] = fifoOut[7][11];
           muxOutConnector[34] = fifoOut[8][11];
           muxOutConnector[35] = fifoOut[9][11];
           muxOutConnector[36] = fifoOut[10][11];
           muxOutConnector[37] = fifoOut[11][11];
           muxOutConnector[38] = fifoOut[12][11];
           muxOutConnector[39] = fifoOut[13][11];
           muxOutConnector[40] = fifoOut[14][11];
           muxOutConnector[41] = fifoOut[15][11];
           muxOutConnector[42] = fifoOut[16][11];
           muxOutConnector[43] = fifoOut[17][11];
           muxOutConnector[44] = fifoOut[18][11];
           muxOutConnector[45] = fifoOut[19][11];
           muxOutConnector[46] = fifoOut[20][11];
           muxOutConnector[47] = fifoOut[21][11];
           muxOutConnector[48] = fifoOut[22][11];
           muxOutConnector[49] = fifoOut[23][11];
           muxOutConnector[50] = fifoOut[24][11];
           muxOutConnector[51] = fifoOut[25][11];
      end
      6: begin
           muxOutConnector[0] = fifoOut[10][0];
           muxOutConnector[1] = fifoOut[11][0];
           muxOutConnector[2] = fifoOut[12][0];
           muxOutConnector[3] = fifoOut[13][0];
           muxOutConnector[4] = fifoOut[14][0];
           muxOutConnector[5] = fifoOut[15][0];
           muxOutConnector[6] = fifoOut[16][0];
           muxOutConnector[7] = fifoOut[17][0];
           muxOutConnector[8] = fifoOut[18][0];
           muxOutConnector[9] = fifoOut[19][0];
           muxOutConnector[10] = fifoOut[20][0];
           muxOutConnector[11] = fifoOut[21][0];
           muxOutConnector[12] = fifoOut[22][0];
           muxOutConnector[13] = fifoOut[23][0];
           muxOutConnector[14] = fifoOut[24][0];
           muxOutConnector[15] = fifoOut[25][0];
           muxOutConnector[16] = fifoOut[26][0];
           muxOutConnector[17] = fifoOut[27][0];
           muxOutConnector[18] = fifoOut[28][0];
           muxOutConnector[19] = fifoOut[29][0];
           muxOutConnector[20] = fifoOut[30][0];
           muxOutConnector[21] = fifoOut[31][0];
           muxOutConnector[22] = fifoOut[0][16];
           muxOutConnector[23] = fifoOut[1][16];
           muxOutConnector[24] = fifoOut[2][16];
           muxOutConnector[25] = fifoOut[3][16];
           muxOutConnector[26] = fifoOut[26][12];
           muxOutConnector[27] = fifoOut[27][12];
           muxOutConnector[28] = fifoOut[28][12];
           muxOutConnector[29] = fifoOut[29][12];
           muxOutConnector[30] = fifoOut[30][12];
           muxOutConnector[31] = fifoOut[31][12];
           muxOutConnector[32] = fifoOut[0][11];
           muxOutConnector[33] = fifoOut[1][11];
           muxOutConnector[34] = fifoOut[2][11];
           muxOutConnector[35] = fifoOut[3][11];
           muxOutConnector[36] = fifoOut[4][11];
           muxOutConnector[37] = fifoOut[5][11];
           muxOutConnector[38] = fifoOut[6][11];
           muxOutConnector[39] = fifoOut[7][11];
           muxOutConnector[40] = fifoOut[8][11];
           muxOutConnector[41] = fifoOut[9][11];
           muxOutConnector[42] = fifoOut[10][11];
           muxOutConnector[43] = fifoOut[11][11];
           muxOutConnector[44] = fifoOut[12][11];
           muxOutConnector[45] = fifoOut[13][11];
           muxOutConnector[46] = fifoOut[14][11];
           muxOutConnector[47] = fifoOut[15][11];
           muxOutConnector[48] = fifoOut[16][11];
           muxOutConnector[49] = fifoOut[17][11];
           muxOutConnector[50] = fifoOut[18][11];
           muxOutConnector[51] = fifoOut[19][11];
      end
      7: begin
           muxOutConnector[0] = fifoOut[4][0];
           muxOutConnector[1] = fifoOut[5][0];
           muxOutConnector[2] = fifoOut[6][0];
           muxOutConnector[3] = fifoOut[7][0];
           muxOutConnector[4] = fifoOut[8][0];
           muxOutConnector[5] = fifoOut[9][0];
           muxOutConnector[6] = fifoOut[10][0];
           muxOutConnector[7] = fifoOut[11][0];
           muxOutConnector[8] = fifoOut[12][0];
           muxOutConnector[9] = fifoOut[13][0];
           muxOutConnector[10] = fifoOut[14][0];
           muxOutConnector[11] = fifoOut[15][0];
           muxOutConnector[12] = fifoOut[16][0];
           muxOutConnector[13] = fifoOut[17][0];
           muxOutConnector[14] = fifoOut[18][0];
           muxOutConnector[15] = fifoOut[19][0];
           muxOutConnector[16] = fifoOut[20][0];
           muxOutConnector[17] = fifoOut[21][0];
           muxOutConnector[18] = fifoOut[22][0];
           muxOutConnector[19] = fifoOut[23][0];
           muxOutConnector[20] = fifoOut[24][0];
           muxOutConnector[21] = fifoOut[25][0];
           muxOutConnector[22] = fifoOut[26][0];
           muxOutConnector[23] = fifoOut[27][0];
           muxOutConnector[24] = fifoOut[28][0];
           muxOutConnector[25] = fifoOut[29][0];
           muxOutConnector[26] = fifoOut[20][12];
           muxOutConnector[27] = fifoOut[21][12];
           muxOutConnector[28] = fifoOut[22][12];
           muxOutConnector[29] = fifoOut[23][12];
           muxOutConnector[30] = fifoOut[24][12];
           muxOutConnector[31] = fifoOut[25][12];
           muxOutConnector[32] = fifoOut[26][12];
           muxOutConnector[33] = fifoOut[27][12];
           muxOutConnector[34] = fifoOut[28][12];
           muxOutConnector[35] = fifoOut[29][12];
           muxOutConnector[36] = fifoOut[30][12];
           muxOutConnector[37] = fifoOut[31][12];
           muxOutConnector[38] = fifoOut[0][11];
           muxOutConnector[39] = fifoOut[1][11];
           muxOutConnector[40] = fifoOut[2][11];
           muxOutConnector[41] = fifoOut[3][11];
           muxOutConnector[42] = fifoOut[4][11];
           muxOutConnector[43] = fifoOut[5][11];
           muxOutConnector[44] = fifoOut[6][11];
           muxOutConnector[45] = fifoOut[7][11];
           muxOutConnector[46] = fifoOut[8][11];
           muxOutConnector[47] = fifoOut[9][11];
           muxOutConnector[48] = fifoOut[10][11];
           muxOutConnector[49] = fifoOut[11][11];
           muxOutConnector[50] = fifoOut[12][11];
           muxOutConnector[51] = fifoOut[13][11];
      end
      8: begin
           muxOutConnector[0] = fifoOut[30][1];
           muxOutConnector[1] = fifoOut[31][1];
           muxOutConnector[2] = fifoOut[0][0];
           muxOutConnector[3] = fifoOut[1][0];
           muxOutConnector[4] = fifoOut[2][0];
           muxOutConnector[5] = fifoOut[3][0];
           muxOutConnector[6] = fifoOut[4][0];
           muxOutConnector[7] = fifoOut[5][0];
           muxOutConnector[8] = fifoOut[6][0];
           muxOutConnector[9] = fifoOut[7][0];
           muxOutConnector[10] = fifoOut[8][0];
           muxOutConnector[11] = fifoOut[9][0];
           muxOutConnector[12] = fifoOut[10][0];
           muxOutConnector[13] = fifoOut[11][0];
           muxOutConnector[14] = fifoOut[12][0];
           muxOutConnector[15] = fifoOut[13][0];
           muxOutConnector[16] = fifoOut[14][0];
           muxOutConnector[17] = fifoOut[15][0];
           muxOutConnector[18] = fifoOut[16][0];
           muxOutConnector[19] = fifoOut[17][0];
           muxOutConnector[20] = fifoOut[18][0];
           muxOutConnector[21] = fifoOut[19][0];
           muxOutConnector[22] = fifoOut[20][0];
           muxOutConnector[23] = fifoOut[21][0];
           muxOutConnector[24] = fifoOut[22][0];
           muxOutConnector[25] = fifoOut[23][0];
           muxOutConnector[26] = fifoOut[14][12];
           muxOutConnector[27] = fifoOut[15][12];
           muxOutConnector[28] = fifoOut[16][12];
           muxOutConnector[29] = fifoOut[17][12];
           muxOutConnector[30] = fifoOut[18][12];
           muxOutConnector[31] = fifoOut[19][12];
           muxOutConnector[32] = fifoOut[20][12];
           muxOutConnector[33] = fifoOut[21][12];
           muxOutConnector[34] = fifoOut[22][12];
           muxOutConnector[35] = fifoOut[23][12];
           muxOutConnector[36] = fifoOut[24][12];
           muxOutConnector[37] = fifoOut[25][12];
           muxOutConnector[38] = fifoOut[26][12];
           muxOutConnector[39] = fifoOut[27][12];
           muxOutConnector[40] = fifoOut[28][12];
           muxOutConnector[41] = fifoOut[29][12];
           muxOutConnector[42] = fifoOut[30][12];
           muxOutConnector[43] = fifoOut[31][12];
           muxOutConnector[44] = fifoOut[0][11];
           muxOutConnector[45] = fifoOut[1][11];
           muxOutConnector[46] = fifoOut[2][11];
           muxOutConnector[47] = fifoOut[3][11];
           muxOutConnector[48] = fifoOut[4][11];
           muxOutConnector[49] = fifoOut[5][11];
           muxOutConnector[50] = fifoOut[6][11];
           muxOutConnector[51] = fifoOut[7][11];
      end
      9: begin
           muxOutConnector[0] = fifoOut[24][1];
           muxOutConnector[1] = fifoOut[25][1];
           muxOutConnector[2] = fifoOut[26][1];
           muxOutConnector[3] = fifoOut[27][1];
           muxOutConnector[4] = fifoOut[28][1];
           muxOutConnector[5] = fifoOut[29][1];
           muxOutConnector[6] = fifoOut[30][1];
           muxOutConnector[7] = fifoOut[31][1];
           muxOutConnector[8] = fifoOut[0][0];
           muxOutConnector[9] = fifoOut[1][0];
           muxOutConnector[10] = fifoOut[2][0];
           muxOutConnector[11] = fifoOut[3][0];
           muxOutConnector[12] = fifoOut[4][0];
           muxOutConnector[13] = fifoOut[5][0];
           muxOutConnector[14] = fifoOut[6][0];
           muxOutConnector[15] = fifoOut[7][0];
           muxOutConnector[16] = fifoOut[8][0];
           muxOutConnector[17] = fifoOut[9][0];
           muxOutConnector[18] = fifoOut[10][0];
           muxOutConnector[19] = fifoOut[11][0];
           muxOutConnector[20] = fifoOut[12][0];
           muxOutConnector[21] = fifoOut[13][0];
           muxOutConnector[22] = fifoOut[14][0];
           muxOutConnector[23] = fifoOut[15][0];
           muxOutConnector[24] = fifoOut[16][0];
           muxOutConnector[25] = fifoOut[17][0];
           muxOutConnector[26] = fifoOut[8][12];
           muxOutConnector[27] = fifoOut[9][12];
           muxOutConnector[28] = fifoOut[10][12];
           muxOutConnector[29] = fifoOut[11][12];
           muxOutConnector[30] = fifoOut[12][12];
           muxOutConnector[31] = fifoOut[13][12];
           muxOutConnector[32] = fifoOut[14][12];
           muxOutConnector[33] = fifoOut[15][12];
           muxOutConnector[34] = fifoOut[16][12];
           muxOutConnector[35] = fifoOut[17][12];
           muxOutConnector[36] = fifoOut[18][12];
           muxOutConnector[37] = fifoOut[19][12];
           muxOutConnector[38] = fifoOut[20][12];
           muxOutConnector[39] = fifoOut[21][12];
           muxOutConnector[40] = fifoOut[22][12];
           muxOutConnector[41] = fifoOut[23][12];
           muxOutConnector[42] = fifoOut[24][12];
           muxOutConnector[43] = fifoOut[25][12];
           muxOutConnector[44] = fifoOut[26][12];
           muxOutConnector[45] = fifoOut[27][12];
           muxOutConnector[46] = fifoOut[28][12];
           muxOutConnector[47] = fifoOut[29][12];
           muxOutConnector[48] = fifoOut[30][12];
           muxOutConnector[49] = fifoOut[31][12];
           muxOutConnector[50] = fifoOut[0][11];
           muxOutConnector[51] = fifoOut[1][11];
      end
      10: begin
           muxOutConnector[0] = fifoOut[18][1];
           muxOutConnector[1] = fifoOut[19][1];
           muxOutConnector[2] = fifoOut[20][1];
           muxOutConnector[3] = fifoOut[21][1];
           muxOutConnector[4] = fifoOut[22][1];
           muxOutConnector[5] = fifoOut[23][1];
           muxOutConnector[6] = fifoOut[24][1];
           muxOutConnector[7] = fifoOut[25][1];
           muxOutConnector[8] = fifoOut[26][1];
           muxOutConnector[9] = fifoOut[27][1];
           muxOutConnector[10] = fifoOut[28][1];
           muxOutConnector[11] = fifoOut[29][1];
           muxOutConnector[12] = fifoOut[30][1];
           muxOutConnector[13] = fifoOut[31][1];
           muxOutConnector[14] = fifoOut[0][0];
           muxOutConnector[15] = fifoOut[1][0];
           muxOutConnector[16] = fifoOut[2][0];
           muxOutConnector[17] = fifoOut[3][0];
           muxOutConnector[18] = fifoOut[4][0];
           muxOutConnector[19] = fifoOut[5][0];
           muxOutConnector[20] = fifoOut[6][0];
           muxOutConnector[21] = fifoOut[7][0];
           muxOutConnector[22] = fifoOut[8][0];
           muxOutConnector[23] = fifoOut[9][0];
           muxOutConnector[24] = fifoOut[10][0];
           muxOutConnector[25] = fifoOut[11][0];
           muxOutConnector[26] = fifoOut[2][12];
           muxOutConnector[27] = fifoOut[3][12];
           muxOutConnector[28] = fifoOut[4][12];
           muxOutConnector[29] = fifoOut[5][12];
           muxOutConnector[30] = fifoOut[6][12];
           muxOutConnector[31] = fifoOut[7][12];
           muxOutConnector[32] = fifoOut[8][12];
           muxOutConnector[33] = fifoOut[9][12];
           muxOutConnector[34] = fifoOut[10][12];
           muxOutConnector[35] = fifoOut[11][12];
           muxOutConnector[36] = fifoOut[12][12];
           muxOutConnector[37] = fifoOut[13][12];
           muxOutConnector[38] = fifoOut[14][12];
           muxOutConnector[39] = fifoOut[15][12];
           muxOutConnector[40] = fifoOut[16][12];
           muxOutConnector[41] = fifoOut[17][12];
           muxOutConnector[42] = fifoOut[18][12];
           muxOutConnector[43] = fifoOut[19][12];
           muxOutConnector[44] = fifoOut[20][12];
           muxOutConnector[45] = fifoOut[21][12];
           muxOutConnector[46] = fifoOut[22][12];
           muxOutConnector[47] = fifoOut[23][12];
           muxOutConnector[48] = fifoOut[24][12];
           muxOutConnector[49] = fifoOut[25][12];
           muxOutConnector[50] = fifoOut[26][12];
           muxOutConnector[51] = fifoOut[27][12];
      end
      11: begin
           muxOutConnector[0] = fifoOut[12][1];
           muxOutConnector[1] = fifoOut[13][1];
           muxOutConnector[2] = fifoOut[14][1];
           muxOutConnector[3] = fifoOut[15][1];
           muxOutConnector[4] = fifoOut[16][1];
           muxOutConnector[5] = fifoOut[17][1];
           muxOutConnector[6] = fifoOut[18][1];
           muxOutConnector[7] = fifoOut[19][1];
           muxOutConnector[8] = fifoOut[20][1];
           muxOutConnector[9] = fifoOut[21][1];
           muxOutConnector[10] = fifoOut[22][1];
           muxOutConnector[11] = fifoOut[23][1];
           muxOutConnector[12] = fifoOut[24][1];
           muxOutConnector[13] = fifoOut[25][1];
           muxOutConnector[14] = fifoOut[26][1];
           muxOutConnector[15] = fifoOut[27][1];
           muxOutConnector[16] = fifoOut[28][1];
           muxOutConnector[17] = fifoOut[29][1];
           muxOutConnector[18] = fifoOut[30][1];
           muxOutConnector[19] = fifoOut[31][1];
           muxOutConnector[20] = fifoOut[0][0];
           muxOutConnector[21] = fifoOut[1][0];
           muxOutConnector[22] = fifoOut[2][0];
           muxOutConnector[23] = fifoOut[3][0];
           muxOutConnector[24] = fifoOut[4][0];
           muxOutConnector[25] = fifoOut[5][0];
           muxOutConnector[26] = fifoOut[28][13];
           muxOutConnector[27] = fifoOut[29][13];
           muxOutConnector[28] = fifoOut[30][13];
           muxOutConnector[29] = fifoOut[31][13];
           muxOutConnector[30] = fifoOut[0][12];
           muxOutConnector[31] = fifoOut[1][12];
           muxOutConnector[32] = fifoOut[2][12];
           muxOutConnector[33] = fifoOut[3][12];
           muxOutConnector[34] = fifoOut[4][12];
           muxOutConnector[35] = fifoOut[5][12];
           muxOutConnector[36] = fifoOut[6][12];
           muxOutConnector[37] = fifoOut[7][12];
           muxOutConnector[38] = fifoOut[8][12];
           muxOutConnector[39] = fifoOut[9][12];
           muxOutConnector[40] = fifoOut[10][12];
           muxOutConnector[41] = fifoOut[11][12];
           muxOutConnector[42] = fifoOut[12][12];
           muxOutConnector[43] = fifoOut[13][12];
           muxOutConnector[44] = fifoOut[14][12];
           muxOutConnector[45] = fifoOut[15][12];
           muxOutConnector[46] = fifoOut[16][12];
           muxOutConnector[47] = fifoOut[17][12];
           muxOutConnector[48] = fifoOut[18][12];
           muxOutConnector[49] = fifoOut[19][12];
           muxOutConnector[50] = fifoOut[20][12];
           muxOutConnector[51] = fifoOut[21][12];
      end
      12: begin
           muxOutConnector[0] = fifoOut[6][1];
           muxOutConnector[1] = fifoOut[7][1];
           muxOutConnector[2] = fifoOut[8][1];
           muxOutConnector[3] = fifoOut[9][1];
           muxOutConnector[4] = fifoOut[10][1];
           muxOutConnector[5] = fifoOut[11][1];
           muxOutConnector[6] = fifoOut[12][1];
           muxOutConnector[7] = fifoOut[13][1];
           muxOutConnector[8] = fifoOut[14][1];
           muxOutConnector[9] = fifoOut[15][1];
           muxOutConnector[10] = fifoOut[16][1];
           muxOutConnector[11] = fifoOut[17][1];
           muxOutConnector[12] = fifoOut[18][1];
           muxOutConnector[13] = fifoOut[19][1];
           muxOutConnector[14] = fifoOut[20][1];
           muxOutConnector[15] = fifoOut[21][1];
           muxOutConnector[16] = fifoOut[22][1];
           muxOutConnector[17] = fifoOut[23][1];
           muxOutConnector[18] = fifoOut[24][1];
           muxOutConnector[19] = fifoOut[25][1];
           muxOutConnector[20] = fifoOut[26][1];
           muxOutConnector[21] = fifoOut[27][1];
           muxOutConnector[22] = fifoOut[28][1];
           muxOutConnector[23] = fifoOut[29][1];
           muxOutConnector[24] = fifoOut[30][1];
           muxOutConnector[25] = fifoOut[31][1];
           muxOutConnector[26] = fifoOut[22][13];
           muxOutConnector[27] = fifoOut[23][13];
           muxOutConnector[28] = fifoOut[24][13];
           muxOutConnector[29] = fifoOut[25][13];
           muxOutConnector[30] = fifoOut[26][13];
           muxOutConnector[31] = fifoOut[27][13];
           muxOutConnector[32] = fifoOut[28][13];
           muxOutConnector[33] = fifoOut[29][13];
           muxOutConnector[34] = fifoOut[30][13];
           muxOutConnector[35] = fifoOut[31][13];
           muxOutConnector[36] = fifoOut[0][12];
           muxOutConnector[37] = fifoOut[1][12];
           muxOutConnector[38] = fifoOut[2][12];
           muxOutConnector[39] = fifoOut[3][12];
           muxOutConnector[40] = fifoOut[4][12];
           muxOutConnector[41] = fifoOut[5][12];
           muxOutConnector[42] = fifoOut[6][12];
           muxOutConnector[43] = fifoOut[7][12];
           muxOutConnector[44] = fifoOut[8][12];
           muxOutConnector[45] = fifoOut[9][12];
           muxOutConnector[46] = fifoOut[10][12];
           muxOutConnector[47] = fifoOut[11][12];
           muxOutConnector[48] = fifoOut[12][12];
           muxOutConnector[49] = maxVal;
           muxOutConnector[50] = maxVal;
           muxOutConnector[51] = maxVal;
      end
      13: begin
           muxOutConnector[0] = fifoOut[0][1];
           muxOutConnector[1] = fifoOut[1][1];
           muxOutConnector[2] = fifoOut[2][1];
           muxOutConnector[3] = fifoOut[3][1];
           muxOutConnector[4] = fifoOut[4][1];
           muxOutConnector[5] = fifoOut[5][1];
           muxOutConnector[6] = fifoOut[6][1];
           muxOutConnector[7] = fifoOut[7][1];
           muxOutConnector[8] = fifoOut[8][1];
           muxOutConnector[9] = fifoOut[9][1];
           muxOutConnector[10] = fifoOut[10][1];
           muxOutConnector[11] = fifoOut[11][1];
           muxOutConnector[12] = fifoOut[12][1];
           muxOutConnector[13] = fifoOut[13][1];
           muxOutConnector[14] = fifoOut[14][1];
           muxOutConnector[15] = fifoOut[15][1];
           muxOutConnector[16] = fifoOut[16][1];
           muxOutConnector[17] = fifoOut[17][1];
           muxOutConnector[18] = fifoOut[18][1];
           muxOutConnector[19] = fifoOut[19][1];
           muxOutConnector[20] = fifoOut[20][1];
           muxOutConnector[21] = fifoOut[21][1];
           muxOutConnector[22] = fifoOut[22][1];
           muxOutConnector[23] = fifoOut[23][1];
           muxOutConnector[24] = fifoOut[24][1];
           muxOutConnector[25] = fifoOut[25][1];
           muxOutConnector[26] = maxVal;
           muxOutConnector[27] = maxVal;
           muxOutConnector[28] = maxVal;
           muxOutConnector[29] = maxVal;
           muxOutConnector[30] = maxVal;
           muxOutConnector[31] = maxVal;
           muxOutConnector[32] = maxVal;
           muxOutConnector[33] = maxVal;
           muxOutConnector[34] = maxVal;
           muxOutConnector[35] = maxVal;
           muxOutConnector[36] = maxVal;
           muxOutConnector[37] = maxVal;
           muxOutConnector[38] = maxVal;
           muxOutConnector[39] = maxVal;
           muxOutConnector[40] = maxVal;
           muxOutConnector[41] = fifoOut[0][11];
           muxOutConnector[42] = fifoOut[1][11];
           muxOutConnector[43] = fifoOut[2][11];
           muxOutConnector[44] = fifoOut[3][11];
           muxOutConnector[45] = fifoOut[4][11];
           muxOutConnector[46] = fifoOut[5][11];
           muxOutConnector[47] = fifoOut[6][11];
           muxOutConnector[48] = fifoOut[7][11];
           muxOutConnector[49] = fifoOut[8][11];
           muxOutConnector[50] = fifoOut[9][11];
           muxOutConnector[51] = fifoOut[10][11];
      end
      14: begin
           muxOutConnector[0] = fifoOut[26][2];
           muxOutConnector[1] = fifoOut[27][2];
           muxOutConnector[2] = fifoOut[28][2];
           muxOutConnector[3] = fifoOut[29][2];
           muxOutConnector[4] = fifoOut[30][2];
           muxOutConnector[5] = fifoOut[31][2];
           muxOutConnector[6] = fifoOut[0][1];
           muxOutConnector[7] = fifoOut[1][1];
           muxOutConnector[8] = fifoOut[2][1];
           muxOutConnector[9] = fifoOut[3][1];
           muxOutConnector[10] = fifoOut[4][1];
           muxOutConnector[11] = fifoOut[5][1];
           muxOutConnector[12] = fifoOut[6][1];
           muxOutConnector[13] = fifoOut[7][1];
           muxOutConnector[14] = fifoOut[8][1];
           muxOutConnector[15] = fifoOut[9][1];
           muxOutConnector[16] = fifoOut[10][1];
           muxOutConnector[17] = fifoOut[11][1];
           muxOutConnector[18] = fifoOut[12][1];
           muxOutConnector[19] = fifoOut[13][1];
           muxOutConnector[20] = fifoOut[14][1];
           muxOutConnector[21] = fifoOut[15][1];
           muxOutConnector[22] = fifoOut[16][1];
           muxOutConnector[23] = fifoOut[17][1];
           muxOutConnector[24] = fifoOut[18][1];
           muxOutConnector[25] = fifoOut[19][1];
           muxOutConnector[26] = fifoOut[11][12];
           muxOutConnector[27] = fifoOut[12][12];
           muxOutConnector[28] = fifoOut[13][12];
           muxOutConnector[29] = fifoOut[14][12];
           muxOutConnector[30] = fifoOut[15][12];
           muxOutConnector[31] = fifoOut[16][12];
           muxOutConnector[32] = fifoOut[17][12];
           muxOutConnector[33] = fifoOut[18][12];
           muxOutConnector[34] = fifoOut[19][12];
           muxOutConnector[35] = fifoOut[20][12];
           muxOutConnector[36] = fifoOut[21][12];
           muxOutConnector[37] = fifoOut[22][12];
           muxOutConnector[38] = fifoOut[23][12];
           muxOutConnector[39] = fifoOut[24][12];
           muxOutConnector[40] = fifoOut[25][12];
           muxOutConnector[41] = fifoOut[26][12];
           muxOutConnector[42] = fifoOut[27][12];
           muxOutConnector[43] = fifoOut[28][12];
           muxOutConnector[44] = fifoOut[29][12];
           muxOutConnector[45] = fifoOut[30][12];
           muxOutConnector[46] = fifoOut[31][12];
           muxOutConnector[47] = fifoOut[0][11];
           muxOutConnector[48] = fifoOut[1][11];
           muxOutConnector[49] = fifoOut[2][11];
           muxOutConnector[50] = fifoOut[3][11];
           muxOutConnector[51] = fifoOut[4][11];
      end
      15: begin
           muxOutConnector[0] = fifoOut[20][2];
           muxOutConnector[1] = fifoOut[21][2];
           muxOutConnector[2] = fifoOut[22][2];
           muxOutConnector[3] = fifoOut[23][2];
           muxOutConnector[4] = fifoOut[24][2];
           muxOutConnector[5] = fifoOut[25][2];
           muxOutConnector[6] = fifoOut[26][2];
           muxOutConnector[7] = fifoOut[27][2];
           muxOutConnector[8] = fifoOut[28][2];
           muxOutConnector[9] = fifoOut[29][2];
           muxOutConnector[10] = fifoOut[30][2];
           muxOutConnector[11] = fifoOut[31][2];
           muxOutConnector[12] = fifoOut[0][1];
           muxOutConnector[13] = fifoOut[1][1];
           muxOutConnector[14] = fifoOut[2][1];
           muxOutConnector[15] = fifoOut[3][1];
           muxOutConnector[16] = fifoOut[4][1];
           muxOutConnector[17] = fifoOut[5][1];
           muxOutConnector[18] = fifoOut[6][1];
           muxOutConnector[19] = fifoOut[7][1];
           muxOutConnector[20] = fifoOut[8][1];
           muxOutConnector[21] = fifoOut[9][1];
           muxOutConnector[22] = fifoOut[10][1];
           muxOutConnector[23] = fifoOut[11][1];
           muxOutConnector[24] = fifoOut[12][1];
           muxOutConnector[25] = fifoOut[13][1];
           muxOutConnector[26] = fifoOut[5][12];
           muxOutConnector[27] = fifoOut[6][12];
           muxOutConnector[28] = fifoOut[7][12];
           muxOutConnector[29] = fifoOut[8][12];
           muxOutConnector[30] = fifoOut[9][12];
           muxOutConnector[31] = fifoOut[10][12];
           muxOutConnector[32] = fifoOut[11][12];
           muxOutConnector[33] = fifoOut[12][12];
           muxOutConnector[34] = fifoOut[13][12];
           muxOutConnector[35] = fifoOut[14][12];
           muxOutConnector[36] = fifoOut[15][12];
           muxOutConnector[37] = fifoOut[16][12];
           muxOutConnector[38] = fifoOut[17][12];
           muxOutConnector[39] = fifoOut[18][12];
           muxOutConnector[40] = fifoOut[19][12];
           muxOutConnector[41] = fifoOut[20][12];
           muxOutConnector[42] = fifoOut[21][12];
           muxOutConnector[43] = fifoOut[22][12];
           muxOutConnector[44] = fifoOut[23][12];
           muxOutConnector[45] = fifoOut[24][12];
           muxOutConnector[46] = fifoOut[25][12];
           muxOutConnector[47] = fifoOut[26][12];
           muxOutConnector[48] = fifoOut[27][12];
           muxOutConnector[49] = fifoOut[28][12];
           muxOutConnector[50] = fifoOut[29][12];
           muxOutConnector[51] = fifoOut[30][12];
      end
      16: begin
           muxOutConnector[0] = fifoOut[14][2];
           muxOutConnector[1] = fifoOut[15][2];
           muxOutConnector[2] = fifoOut[16][2];
           muxOutConnector[3] = fifoOut[17][2];
           muxOutConnector[4] = fifoOut[18][2];
           muxOutConnector[5] = fifoOut[19][2];
           muxOutConnector[6] = fifoOut[20][2];
           muxOutConnector[7] = fifoOut[21][2];
           muxOutConnector[8] = fifoOut[22][2];
           muxOutConnector[9] = fifoOut[23][2];
           muxOutConnector[10] = fifoOut[24][2];
           muxOutConnector[11] = fifoOut[25][2];
           muxOutConnector[12] = fifoOut[26][2];
           muxOutConnector[13] = fifoOut[27][2];
           muxOutConnector[14] = fifoOut[28][2];
           muxOutConnector[15] = fifoOut[29][2];
           muxOutConnector[16] = fifoOut[30][2];
           muxOutConnector[17] = fifoOut[31][2];
           muxOutConnector[18] = fifoOut[0][1];
           muxOutConnector[19] = fifoOut[1][1];
           muxOutConnector[20] = fifoOut[2][1];
           muxOutConnector[21] = fifoOut[3][1];
           muxOutConnector[22] = fifoOut[4][1];
           muxOutConnector[23] = fifoOut[5][1];
           muxOutConnector[24] = fifoOut[6][1];
           muxOutConnector[25] = fifoOut[7][1];
           muxOutConnector[26] = fifoOut[31][13];
           muxOutConnector[27] = fifoOut[0][12];
           muxOutConnector[28] = fifoOut[1][12];
           muxOutConnector[29] = fifoOut[2][12];
           muxOutConnector[30] = fifoOut[3][12];
           muxOutConnector[31] = fifoOut[4][12];
           muxOutConnector[32] = fifoOut[5][12];
           muxOutConnector[33] = fifoOut[6][12];
           muxOutConnector[34] = fifoOut[7][12];
           muxOutConnector[35] = fifoOut[8][12];
           muxOutConnector[36] = fifoOut[9][12];
           muxOutConnector[37] = fifoOut[10][12];
           muxOutConnector[38] = fifoOut[11][12];
           muxOutConnector[39] = fifoOut[12][12];
           muxOutConnector[40] = fifoOut[13][12];
           muxOutConnector[41] = fifoOut[14][12];
           muxOutConnector[42] = fifoOut[15][12];
           muxOutConnector[43] = fifoOut[16][12];
           muxOutConnector[44] = fifoOut[17][12];
           muxOutConnector[45] = fifoOut[18][12];
           muxOutConnector[46] = fifoOut[19][12];
           muxOutConnector[47] = fifoOut[20][12];
           muxOutConnector[48] = fifoOut[21][12];
           muxOutConnector[49] = fifoOut[22][12];
           muxOutConnector[50] = fifoOut[23][12];
           muxOutConnector[51] = fifoOut[24][12];
      end
      17: begin
           muxOutConnector[0] = fifoOut[8][2];
           muxOutConnector[1] = fifoOut[9][2];
           muxOutConnector[2] = fifoOut[10][2];
           muxOutConnector[3] = fifoOut[11][2];
           muxOutConnector[4] = fifoOut[12][2];
           muxOutConnector[5] = fifoOut[13][2];
           muxOutConnector[6] = fifoOut[14][2];
           muxOutConnector[7] = fifoOut[15][2];
           muxOutConnector[8] = fifoOut[16][2];
           muxOutConnector[9] = fifoOut[17][2];
           muxOutConnector[10] = fifoOut[18][2];
           muxOutConnector[11] = fifoOut[19][2];
           muxOutConnector[12] = fifoOut[20][2];
           muxOutConnector[13] = fifoOut[21][2];
           muxOutConnector[14] = fifoOut[22][2];
           muxOutConnector[15] = fifoOut[23][2];
           muxOutConnector[16] = fifoOut[24][2];
           muxOutConnector[17] = fifoOut[25][2];
           muxOutConnector[18] = fifoOut[26][2];
           muxOutConnector[19] = fifoOut[27][2];
           muxOutConnector[20] = fifoOut[28][2];
           muxOutConnector[21] = fifoOut[29][2];
           muxOutConnector[22] = fifoOut[30][2];
           muxOutConnector[23] = fifoOut[31][2];
           muxOutConnector[24] = fifoOut[0][1];
           muxOutConnector[25] = fifoOut[1][1];
           muxOutConnector[26] = fifoOut[25][13];
           muxOutConnector[27] = fifoOut[26][13];
           muxOutConnector[28] = fifoOut[27][13];
           muxOutConnector[29] = fifoOut[28][13];
           muxOutConnector[30] = fifoOut[29][13];
           muxOutConnector[31] = fifoOut[30][13];
           muxOutConnector[32] = fifoOut[31][13];
           muxOutConnector[33] = fifoOut[0][12];
           muxOutConnector[34] = fifoOut[1][12];
           muxOutConnector[35] = fifoOut[2][12];
           muxOutConnector[36] = fifoOut[3][12];
           muxOutConnector[37] = fifoOut[4][12];
           muxOutConnector[38] = fifoOut[5][12];
           muxOutConnector[39] = fifoOut[6][12];
           muxOutConnector[40] = fifoOut[7][12];
           muxOutConnector[41] = fifoOut[8][12];
           muxOutConnector[42] = fifoOut[9][12];
           muxOutConnector[43] = fifoOut[10][12];
           muxOutConnector[44] = fifoOut[11][12];
           muxOutConnector[45] = fifoOut[12][12];
           muxOutConnector[46] = fifoOut[13][12];
           muxOutConnector[47] = fifoOut[14][12];
           muxOutConnector[48] = fifoOut[15][12];
           muxOutConnector[49] = fifoOut[16][12];
           muxOutConnector[50] = fifoOut[17][12];
           muxOutConnector[51] = fifoOut[18][12];
      end
      18: begin
           muxOutConnector[0] = fifoOut[2][2];
           muxOutConnector[1] = fifoOut[3][2];
           muxOutConnector[2] = fifoOut[4][2];
           muxOutConnector[3] = fifoOut[5][2];
           muxOutConnector[4] = fifoOut[6][2];
           muxOutConnector[5] = fifoOut[7][2];
           muxOutConnector[6] = fifoOut[8][2];
           muxOutConnector[7] = fifoOut[9][2];
           muxOutConnector[8] = fifoOut[10][2];
           muxOutConnector[9] = fifoOut[11][2];
           muxOutConnector[10] = fifoOut[12][2];
           muxOutConnector[11] = fifoOut[13][2];
           muxOutConnector[12] = fifoOut[14][2];
           muxOutConnector[13] = fifoOut[15][2];
           muxOutConnector[14] = fifoOut[16][2];
           muxOutConnector[15] = fifoOut[17][2];
           muxOutConnector[16] = fifoOut[18][2];
           muxOutConnector[17] = fifoOut[19][2];
           muxOutConnector[18] = fifoOut[20][2];
           muxOutConnector[19] = fifoOut[21][2];
           muxOutConnector[20] = fifoOut[22][2];
           muxOutConnector[21] = fifoOut[23][2];
           muxOutConnector[22] = fifoOut[24][2];
           muxOutConnector[23] = fifoOut[25][2];
           muxOutConnector[24] = fifoOut[26][2];
           muxOutConnector[25] = fifoOut[27][2];
           muxOutConnector[26] = fifoOut[19][13];
           muxOutConnector[27] = fifoOut[20][13];
           muxOutConnector[28] = fifoOut[21][13];
           muxOutConnector[29] = fifoOut[22][13];
           muxOutConnector[30] = fifoOut[23][13];
           muxOutConnector[31] = fifoOut[24][13];
           muxOutConnector[32] = fifoOut[25][13];
           muxOutConnector[33] = fifoOut[26][13];
           muxOutConnector[34] = fifoOut[27][13];
           muxOutConnector[35] = fifoOut[28][13];
           muxOutConnector[36] = fifoOut[29][13];
           muxOutConnector[37] = fifoOut[30][13];
           muxOutConnector[38] = fifoOut[31][13];
           muxOutConnector[39] = fifoOut[0][12];
           muxOutConnector[40] = fifoOut[1][12];
           muxOutConnector[41] = fifoOut[2][12];
           muxOutConnector[42] = fifoOut[3][12];
           muxOutConnector[43] = fifoOut[4][12];
           muxOutConnector[44] = fifoOut[5][12];
           muxOutConnector[45] = fifoOut[6][12];
           muxOutConnector[46] = fifoOut[7][12];
           muxOutConnector[47] = fifoOut[8][12];
           muxOutConnector[48] = fifoOut[9][12];
           muxOutConnector[49] = fifoOut[10][12];
           muxOutConnector[50] = fifoOut[11][12];
           muxOutConnector[51] = fifoOut[12][12];
      end
      19: begin
           muxOutConnector[0] = fifoOut[28][3];
           muxOutConnector[1] = fifoOut[29][3];
           muxOutConnector[2] = fifoOut[30][3];
           muxOutConnector[3] = fifoOut[31][3];
           muxOutConnector[4] = fifoOut[0][2];
           muxOutConnector[5] = fifoOut[1][2];
           muxOutConnector[6] = fifoOut[2][2];
           muxOutConnector[7] = fifoOut[3][2];
           muxOutConnector[8] = fifoOut[4][2];
           muxOutConnector[9] = fifoOut[5][2];
           muxOutConnector[10] = fifoOut[6][2];
           muxOutConnector[11] = fifoOut[7][2];
           muxOutConnector[12] = fifoOut[8][2];
           muxOutConnector[13] = fifoOut[9][2];
           muxOutConnector[14] = fifoOut[10][2];
           muxOutConnector[15] = fifoOut[11][2];
           muxOutConnector[16] = fifoOut[12][2];
           muxOutConnector[17] = fifoOut[31][2];
           muxOutConnector[18] = fifoOut[31][2];
           muxOutConnector[19] = fifoOut[31][2];
           muxOutConnector[20] = fifoOut[31][2];
           muxOutConnector[21] = fifoOut[31][2];
           muxOutConnector[22] = fifoOut[31][2];
           muxOutConnector[23] = fifoOut[31][2];
           muxOutConnector[24] = fifoOut[31][2];
           muxOutConnector[25] = fifoOut[31][2];
           muxOutConnector[26] = fifoOut[13][13];
           muxOutConnector[27] = fifoOut[14][13];
           muxOutConnector[28] = fifoOut[15][13];
           muxOutConnector[29] = fifoOut[16][13];
           muxOutConnector[30] = fifoOut[17][13];
           muxOutConnector[31] = fifoOut[18][13];
           muxOutConnector[32] = fifoOut[19][13];
           muxOutConnector[33] = fifoOut[20][13];
           muxOutConnector[34] = fifoOut[21][13];
           muxOutConnector[35] = fifoOut[22][13];
           muxOutConnector[36] = fifoOut[23][13];
           muxOutConnector[37] = fifoOut[24][13];
           muxOutConnector[38] = fifoOut[25][13];
           muxOutConnector[39] = fifoOut[26][13];
           muxOutConnector[40] = fifoOut[27][13];
           muxOutConnector[41] = fifoOut[28][13];
           muxOutConnector[42] = fifoOut[29][13];
           muxOutConnector[43] = fifoOut[31][2];
           muxOutConnector[44] = fifoOut[31][2];
           muxOutConnector[45] = fifoOut[31][2];
           muxOutConnector[46] = fifoOut[31][2];
           muxOutConnector[47] = fifoOut[31][2];
           muxOutConnector[48] = fifoOut[31][2];
           muxOutConnector[49] = fifoOut[31][2];
           muxOutConnector[50] = fifoOut[31][2];
           muxOutConnector[51] = fifoOut[31][2];
      end
      default: begin
            for(i=0;i<muxOutSymbols;i=i+1)begin
             muxOutConnector[i] = 0;
           end
      end
  endcase
 end
      default: begin
            for(i=0;i<muxOutSymbols;i=i+1)begin
             muxOutConnector[i] = 0;
           end
      end
 endcase
end
endmodule
                                                                                                                                  12];
              muxOutConnector[51] = fifoOut[12][12];
         end
         19: begin
              muxOutConnector[0] = fifoOut[28][3];
              muxOutConnector[1] = fifoOut[29][3];
              muxOutConnector[2] = fifoOut[30][3];
              muxOutConnector[3] = fifoOut[31][3];
              muxOutConnector[4] = fifoOut[0][2];
              muxOutConnector[5] = fifoOut[1][2];
              muxOutConnector[6] = fifoOut[2][2];
              muxOutConnector[7] = fifoOut[3][2];
              muxOutConnector[8] = fifoOut[4][2];
              muxOutConnector[9] = fifoOut[5][2];
              muxOutConnector[10] = fifoOut[6][2];
              muxOutConnector[11] = fifoOut[7][2];
              muxOutConnector[12] = fifoOut[8][2];
              muxOutConnector[13] = fifoOut[9][2];
              muxOutConnector[14] = fifoOut[10][2];
              muxOutConnector[15] = fifoOut[11][2];
              muxOutConnector[16] = fifoOut[12][2];
              muxOutConnector[17] = fifoOut[31][2];
              muxOutConnector[18] = fifoOut[31][2];
              muxOutConnector[19] = fifoOut[31][2];
              muxOutConnector[20] = fifoOut[31][2];
              muxOutConnector[21] = fifoOut[31][2];
              muxOutConnector[22] = fifoOut[31][2];
              muxOutConnector[23] = fifoOut[31][2];
              muxOutConnector[24] = fifoOut[31][2];
              muxOutConnector[25] = fifoOut[31][2];
              muxOutConnector[26] = fifoOut[13][13];
              muxOutConnector[27] = fifoOut[14][13];
              muxOutConnector[28] = fifoOut[15][13];
              muxOutConnector[29] = fifoOut[16][13];
              muxOutConnector[30] = fifoOut[17][13];
              muxOutConnector[31] = fifoOut[18][13];
              muxOutConnector[32] = fifoOut[19][13];
              muxOutConnector[33] = fifoOut[20][13];
              muxOutConnector[34] = fifoOut[21][13];
              muxOutConnector[35] = fifoOut[22][13];
              muxOutConnector[36] = fifoOut[23][13];
              muxOutConnector[37] = fifoOut[24][13];
              muxOutConnector[38] = fifoOut[25][13];
              muxOutConnector[39] = fifoOut[26][13];
              muxOutConnector[40] = fifoOut[27][13];
              muxOutConnector[41] = fifoOut[28][13];
              muxOutConnector[42] = fifoOut[29][13];
              muxOutConnector[43] = fifoOut[31][2];
              muxOutConnector[44] = fifoOut[31][2];
              muxOutConnector[45] = fifoOut[31][2];
              muxOutConnector[46] = fifoOut[31][2];
              muxOutConnector[47] = fifoOut[31][2];
              muxOutConnector[48] = fifoOut[31][2];
              muxOutConnector[49] = fifoOut[31][2];
              muxOutConnector[50] = fifoOut[31][2];
              muxOutConnector[51] = fifoOut[31][2];
         end
         default: begin
               for(i=0;i<muxOutSymbols;i=i+1)begin
                muxOutConnector[i] = 0;
              end
         end
     endcase
    end
         default: begin
               for(i=0;i<muxOutSymbols;i=i+1)begin
                muxOutConnector[i] = 0;
              end
         end
    endcase
end
endmodule
