`timescale 1ns / 1ps
module LMem1To0_511_circ9_yesshift_nounload_scripted(
        muxOut,
        ly0In,
        wr_en,
        feedback_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 15;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

input feedback_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        if(feedback_en) begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= fifoOut[i][c-1];
         end
        end
        else begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= ly0InConnector[i];
         end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[43][4];
              muxOutConnector[45] = fifoOut[44][4];
              muxOutConnector[46] = fifoOut[45][4];
              muxOutConnector[47] = fifoOut[46][4];
              muxOutConnector[48] = fifoOut[47][4];
              muxOutConnector[49] = fifoOut[48][4];
              muxOutConnector[50] = fifoOut[49][4];
              muxOutConnector[51] = fifoOut[50][4];
       end
       1: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[43][4];
              muxOutConnector[45] = fifoOut[44][4];
              muxOutConnector[46] = fifoOut[45][4];
              muxOutConnector[47] = fifoOut[46][4];
              muxOutConnector[48] = fifoOut[47][4];
              muxOutConnector[49] = fifoOut[48][4];
              muxOutConnector[50] = fifoOut[49][4];
              muxOutConnector[51] = fifoOut[50][4];
       end
       2: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[43][4];
              muxOutConnector[45] = fifoOut[44][4];
              muxOutConnector[46] = fifoOut[45][4];
              muxOutConnector[47] = fifoOut[46][4];
              muxOutConnector[48] = fifoOut[47][4];
              muxOutConnector[49] = fifoOut[48][4];
              muxOutConnector[50] = fifoOut[49][4];
              muxOutConnector[51] = fifoOut[50][4];
       end
       3: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[43][4];
              muxOutConnector[45] = fifoOut[44][4];
              muxOutConnector[46] = fifoOut[45][4];
              muxOutConnector[47] = fifoOut[46][4];
              muxOutConnector[48] = fifoOut[47][4];
              muxOutConnector[49] = fifoOut[48][4];
              muxOutConnector[50] = fifoOut[49][4];
              muxOutConnector[51] = fifoOut[50][4];
       end
       4: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[51][5];
              muxOutConnector[27] = fifoOut[26][4];
              muxOutConnector[28] = fifoOut[27][4];
              muxOutConnector[29] = fifoOut[28][4];
              muxOutConnector[30] = fifoOut[29][4];
              muxOutConnector[31] = fifoOut[30][4];
              muxOutConnector[32] = fifoOut[31][4];
              muxOutConnector[33] = fifoOut[32][4];
              muxOutConnector[34] = fifoOut[33][4];
              muxOutConnector[35] = fifoOut[34][4];
              muxOutConnector[36] = fifoOut[35][4];
              muxOutConnector[37] = fifoOut[36][4];
              muxOutConnector[38] = fifoOut[37][4];
              muxOutConnector[39] = fifoOut[38][4];
              muxOutConnector[40] = fifoOut[39][4];
              muxOutConnector[41] = fifoOut[40][4];
              muxOutConnector[42] = fifoOut[41][4];
              muxOutConnector[43] = fifoOut[42][4];
              muxOutConnector[44] = fifoOut[19][3];
              muxOutConnector[45] = fifoOut[20][3];
              muxOutConnector[46] = fifoOut[21][3];
              muxOutConnector[47] = fifoOut[22][3];
              muxOutConnector[48] = fifoOut[23][3];
              muxOutConnector[49] = fifoOut[24][3];
              muxOutConnector[50] = fifoOut[25][3];
              muxOutConnector[51] = fifoOut[0][2];
       end
       5: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][3];
              muxOutConnector[27] = fifoOut[2][3];
              muxOutConnector[28] = fifoOut[3][3];
              muxOutConnector[29] = fifoOut[4][3];
              muxOutConnector[30] = fifoOut[5][3];
              muxOutConnector[31] = fifoOut[6][3];
              muxOutConnector[32] = fifoOut[7][3];
              muxOutConnector[33] = fifoOut[8][3];
              muxOutConnector[34] = fifoOut[9][3];
              muxOutConnector[35] = fifoOut[10][3];
              muxOutConnector[36] = fifoOut[11][3];
              muxOutConnector[37] = fifoOut[12][3];
              muxOutConnector[38] = fifoOut[13][3];
              muxOutConnector[39] = fifoOut[14][3];
              muxOutConnector[40] = fifoOut[15][3];
              muxOutConnector[41] = fifoOut[16][3];
              muxOutConnector[42] = fifoOut[17][3];
              muxOutConnector[43] = fifoOut[18][3];
              muxOutConnector[44] = fifoOut[19][3];
              muxOutConnector[45] = fifoOut[20][3];
              muxOutConnector[46] = fifoOut[21][3];
              muxOutConnector[47] = fifoOut[22][3];
              muxOutConnector[48] = fifoOut[23][3];
              muxOutConnector[49] = fifoOut[24][3];
              muxOutConnector[50] = fifoOut[25][3];
              muxOutConnector[51] = fifoOut[0][2];
       end
       6: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][3];
              muxOutConnector[27] = fifoOut[2][3];
              muxOutConnector[28] = fifoOut[3][3];
              muxOutConnector[29] = fifoOut[4][3];
              muxOutConnector[30] = fifoOut[5][3];
              muxOutConnector[31] = fifoOut[6][3];
              muxOutConnector[32] = fifoOut[7][3];
              muxOutConnector[33] = fifoOut[8][3];
              muxOutConnector[34] = fifoOut[9][3];
              muxOutConnector[35] = fifoOut[10][3];
              muxOutConnector[36] = fifoOut[11][3];
              muxOutConnector[37] = fifoOut[12][3];
              muxOutConnector[38] = fifoOut[13][3];
              muxOutConnector[39] = fifoOut[14][3];
              muxOutConnector[40] = fifoOut[15][3];
              muxOutConnector[41] = fifoOut[16][3];
              muxOutConnector[42] = fifoOut[17][3];
              muxOutConnector[43] = fifoOut[18][3];
              muxOutConnector[44] = fifoOut[19][3];
              muxOutConnector[45] = fifoOut[20][3];
              muxOutConnector[46] = fifoOut[21][3];
              muxOutConnector[47] = fifoOut[22][3];
              muxOutConnector[48] = fifoOut[23][3];
              muxOutConnector[49] = fifoOut[24][3];
              muxOutConnector[50] = fifoOut[25][3];
              muxOutConnector[51] = fifoOut[0][2];
       end
       7: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][3];
              muxOutConnector[27] = fifoOut[2][3];
              muxOutConnector[28] = fifoOut[3][3];
              muxOutConnector[29] = fifoOut[4][3];
              muxOutConnector[30] = fifoOut[5][3];
              muxOutConnector[31] = fifoOut[6][3];
              muxOutConnector[32] = fifoOut[7][3];
              muxOutConnector[33] = fifoOut[8][3];
              muxOutConnector[34] = fifoOut[9][3];
              muxOutConnector[35] = fifoOut[10][3];
              muxOutConnector[36] = fifoOut[11][3];
              muxOutConnector[37] = fifoOut[12][3];
              muxOutConnector[38] = fifoOut[13][3];
              muxOutConnector[39] = fifoOut[14][3];
              muxOutConnector[40] = fifoOut[15][3];
              muxOutConnector[41] = fifoOut[16][3];
              muxOutConnector[42] = fifoOut[17][3];
              muxOutConnector[43] = fifoOut[18][3];
              muxOutConnector[44] = fifoOut[19][3];
              muxOutConnector[45] = fifoOut[20][3];
              muxOutConnector[46] = fifoOut[21][3];
              muxOutConnector[47] = fifoOut[22][3];
              muxOutConnector[48] = fifoOut[23][3];
              muxOutConnector[49] = fifoOut[24][3];
              muxOutConnector[50] = fifoOut[25][3];
              muxOutConnector[51] = fifoOut[0][2];
       end
       8: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[17][9];
              muxOutConnector[16] = fifoOut[18][9];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][3];
              muxOutConnector[27] = fifoOut[2][3];
              muxOutConnector[28] = fifoOut[3][3];
              muxOutConnector[29] = fifoOut[4][3];
              muxOutConnector[30] = fifoOut[5][3];
              muxOutConnector[31] = fifoOut[6][3];
              muxOutConnector[32] = fifoOut[7][3];
              muxOutConnector[33] = fifoOut[8][3];
              muxOutConnector[34] = fifoOut[9][3];
              muxOutConnector[35] = fifoOut[10][3];
              muxOutConnector[36] = fifoOut[11][3];
              muxOutConnector[37] = fifoOut[12][3];
              muxOutConnector[38] = fifoOut[13][3];
              muxOutConnector[39] = fifoOut[14][3];
              muxOutConnector[40] = fifoOut[15][3];
              muxOutConnector[41] = fifoOut[16][3];
              muxOutConnector[42] = fifoOut[17][3];
              muxOutConnector[43] = fifoOut[18][3];
              muxOutConnector[44] = fifoOut[19][3];
              muxOutConnector[45] = fifoOut[20][3];
              muxOutConnector[46] = fifoOut[21][3];
              muxOutConnector[47] = fifoOut[22][3];
              muxOutConnector[48] = fifoOut[23][3];
              muxOutConnector[49] = fifoOut[24][3];
              muxOutConnector[50] = fifoOut[25][3];
              muxOutConnector[51] = fifoOut[0][2];
       end
       9: begin
              muxOutConnector[0] = fifoOut[2][9];
              muxOutConnector[1] = fifoOut[3][9];
              muxOutConnector[2] = fifoOut[4][9];
              muxOutConnector[3] = fifoOut[5][9];
              muxOutConnector[4] = fifoOut[6][9];
              muxOutConnector[5] = fifoOut[7][9];
              muxOutConnector[6] = fifoOut[8][9];
              muxOutConnector[7] = fifoOut[9][9];
              muxOutConnector[8] = fifoOut[10][9];
              muxOutConnector[9] = fifoOut[11][9];
              muxOutConnector[10] = fifoOut[12][9];
              muxOutConnector[11] = fifoOut[13][9];
              muxOutConnector[12] = fifoOut[14][9];
              muxOutConnector[13] = fifoOut[15][9];
              muxOutConnector[14] = fifoOut[16][9];
              muxOutConnector[15] = fifoOut[50][0];
              muxOutConnector[16] = fifoOut[51][0];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[1][3];
              muxOutConnector[27] = fifoOut[2][3];
              muxOutConnector[28] = fifoOut[3][3];
              muxOutConnector[29] = fifoOut[4][3];
              muxOutConnector[30] = fifoOut[5][3];
              muxOutConnector[31] = fifoOut[6][3];
              muxOutConnector[32] = fifoOut[7][3];
              muxOutConnector[33] = fifoOut[8][3];
              muxOutConnector[34] = fifoOut[9][3];
              muxOutConnector[35] = fifoOut[10][3];
              muxOutConnector[36] = fifoOut[11][3];
              muxOutConnector[37] = fifoOut[12][3];
              muxOutConnector[38] = fifoOut[13][3];
              muxOutConnector[39] = fifoOut[14][3];
              muxOutConnector[40] = fifoOut[15][3];
              muxOutConnector[41] = fifoOut[16][3];
              muxOutConnector[42] = fifoOut[17][3];
              muxOutConnector[43] = fifoOut[18][3];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       10: begin
              muxOutConnector[0] = fifoOut[35][0];
              muxOutConnector[1] = fifoOut[36][0];
              muxOutConnector[2] = fifoOut[37][0];
              muxOutConnector[3] = fifoOut[38][0];
              muxOutConnector[4] = fifoOut[39][0];
              muxOutConnector[5] = fifoOut[40][0];
              muxOutConnector[6] = fifoOut[41][0];
              muxOutConnector[7] = fifoOut[42][0];
              muxOutConnector[8] = fifoOut[43][0];
              muxOutConnector[9] = fifoOut[44][0];
              muxOutConnector[10] = fifoOut[45][0];
              muxOutConnector[11] = fifoOut[46][0];
              muxOutConnector[12] = fifoOut[47][0];
              muxOutConnector[13] = fifoOut[48][0];
              muxOutConnector[14] = fifoOut[49][0];
              muxOutConnector[15] = fifoOut[50][0];
              muxOutConnector[16] = fifoOut[51][0];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       11: begin
              muxOutConnector[0] = fifoOut[35][0];
              muxOutConnector[1] = fifoOut[36][0];
              muxOutConnector[2] = fifoOut[37][0];
              muxOutConnector[3] = fifoOut[38][0];
              muxOutConnector[4] = fifoOut[39][0];
              muxOutConnector[5] = fifoOut[40][0];
              muxOutConnector[6] = fifoOut[41][0];
              muxOutConnector[7] = fifoOut[42][0];
              muxOutConnector[8] = fifoOut[43][0];
              muxOutConnector[9] = fifoOut[44][0];
              muxOutConnector[10] = fifoOut[45][0];
              muxOutConnector[11] = fifoOut[46][0];
              muxOutConnector[12] = fifoOut[47][0];
              muxOutConnector[13] = fifoOut[48][0];
              muxOutConnector[14] = fifoOut[49][0];
              muxOutConnector[15] = fifoOut[50][0];
              muxOutConnector[16] = fifoOut[51][0];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       12: begin
              muxOutConnector[0] = fifoOut[35][0];
              muxOutConnector[1] = fifoOut[36][0];
              muxOutConnector[2] = fifoOut[37][0];
              muxOutConnector[3] = fifoOut[38][0];
              muxOutConnector[4] = fifoOut[39][0];
              muxOutConnector[5] = fifoOut[40][0];
              muxOutConnector[6] = fifoOut[41][0];
              muxOutConnector[7] = fifoOut[42][0];
              muxOutConnector[8] = fifoOut[43][0];
              muxOutConnector[9] = fifoOut[44][0];
              muxOutConnector[10] = fifoOut[45][0];
              muxOutConnector[11] = fifoOut[46][0];
              muxOutConnector[12] = fifoOut[47][0];
              muxOutConnector[13] = fifoOut[48][0];
              muxOutConnector[14] = fifoOut[49][0];
              muxOutConnector[15] = fifoOut[50][0];
              muxOutConnector[16] = fifoOut[51][0];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       13: begin
              muxOutConnector[0] = fifoOut[35][0];
              muxOutConnector[1] = fifoOut[36][0];
              muxOutConnector[2] = fifoOut[37][0];
              muxOutConnector[3] = fifoOut[38][0];
              muxOutConnector[4] = fifoOut[39][0];
              muxOutConnector[5] = fifoOut[40][0];
              muxOutConnector[6] = fifoOut[41][0];
              muxOutConnector[7] = fifoOut[42][0];
              muxOutConnector[8] = fifoOut[43][0];
              muxOutConnector[9] = fifoOut[44][0];
              muxOutConnector[10] = fifoOut[45][0];
              muxOutConnector[11] = fifoOut[46][0];
              muxOutConnector[12] = fifoOut[47][0];
              muxOutConnector[13] = fifoOut[48][0];
              muxOutConnector[14] = fifoOut[49][0];
              muxOutConnector[15] = fifoOut[50][0];
              muxOutConnector[16] = fifoOut[51][0];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       14: begin
              muxOutConnector[0] = fifoOut[35][0];
              muxOutConnector[1] = fifoOut[36][0];
              muxOutConnector[2] = fifoOut[37][0];
              muxOutConnector[3] = fifoOut[38][0];
              muxOutConnector[4] = fifoOut[39][0];
              muxOutConnector[5] = fifoOut[40][0];
              muxOutConnector[6] = fifoOut[41][0];
              muxOutConnector[7] = fifoOut[42][0];
              muxOutConnector[8] = fifoOut[43][0];
              muxOutConnector[9] = fifoOut[44][0];
              muxOutConnector[10] = fifoOut[45][0];
              muxOutConnector[11] = fifoOut[46][0];
              muxOutConnector[12] = fifoOut[47][0];
              muxOutConnector[13] = fifoOut[48][0];
              muxOutConnector[14] = fifoOut[49][0];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[26][14];
              muxOutConnector[18] = fifoOut[27][14];
              muxOutConnector[19] = fifoOut[28][14];
              muxOutConnector[20] = fifoOut[29][14];
              muxOutConnector[21] = fifoOut[30][14];
              muxOutConnector[22] = fifoOut[31][14];
              muxOutConnector[23] = fifoOut[32][14];
              muxOutConnector[24] = fifoOut[33][14];
              muxOutConnector[25] = fifoOut[34][14];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       15: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[2][13];
              muxOutConnector[18] = fifoOut[3][13];
              muxOutConnector[19] = fifoOut[4][13];
              muxOutConnector[20] = fifoOut[5][13];
              muxOutConnector[21] = fifoOut[6][13];
              muxOutConnector[22] = fifoOut[7][13];
              muxOutConnector[23] = fifoOut[8][13];
              muxOutConnector[24] = fifoOut[9][13];
              muxOutConnector[25] = fifoOut[10][13];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       16: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[2][13];
              muxOutConnector[18] = fifoOut[3][13];
              muxOutConnector[19] = fifoOut[4][13];
              muxOutConnector[20] = fifoOut[5][13];
              muxOutConnector[21] = fifoOut[6][13];
              muxOutConnector[22] = fifoOut[7][13];
              muxOutConnector[23] = fifoOut[8][13];
              muxOutConnector[24] = fifoOut[9][13];
              muxOutConnector[25] = fifoOut[10][13];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       17: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[2][13];
              muxOutConnector[18] = fifoOut[3][13];
              muxOutConnector[19] = fifoOut[4][13];
              muxOutConnector[20] = fifoOut[5][13];
              muxOutConnector[21] = fifoOut[6][13];
              muxOutConnector[22] = fifoOut[7][13];
              muxOutConnector[23] = fifoOut[8][13];
              muxOutConnector[24] = fifoOut[9][13];
              muxOutConnector[25] = fifoOut[10][13];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       18: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = fifoOut[2][13];
              muxOutConnector[18] = fifoOut[3][13];
              muxOutConnector[19] = fifoOut[4][13];
              muxOutConnector[20] = fifoOut[5][13];
              muxOutConnector[21] = fifoOut[6][13];
              muxOutConnector[22] = fifoOut[7][13];
              muxOutConnector[23] = fifoOut[8][13];
              muxOutConnector[24] = fifoOut[9][13];
              muxOutConnector[25] = fifoOut[10][13];
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = fifoOut[51][9];
              muxOutConnector[44] = fifoOut[26][8];
              muxOutConnector[45] = fifoOut[27][8];
              muxOutConnector[46] = fifoOut[28][8];
              muxOutConnector[47] = fifoOut[29][8];
              muxOutConnector[48] = fifoOut[30][8];
              muxOutConnector[49] = fifoOut[31][8];
              muxOutConnector[50] = fifoOut[32][8];
              muxOutConnector[51] = fifoOut[33][8];
       end
       19: begin
              muxOutConnector[0] = fifoOut[11][14];
              muxOutConnector[1] = fifoOut[12][14];
              muxOutConnector[2] = fifoOut[13][14];
              muxOutConnector[3] = fifoOut[14][14];
              muxOutConnector[4] = fifoOut[15][14];
              muxOutConnector[5] = fifoOut[16][14];
              muxOutConnector[6] = fifoOut[17][14];
              muxOutConnector[7] = fifoOut[18][14];
              muxOutConnector[8] = fifoOut[19][14];
              muxOutConnector[9] = fifoOut[20][14];
              muxOutConnector[10] = fifoOut[21][14];
              muxOutConnector[11] = fifoOut[22][14];
              muxOutConnector[12] = fifoOut[23][14];
              muxOutConnector[13] = fifoOut[24][14];
              muxOutConnector[14] = fifoOut[25][14];
              muxOutConnector[15] = fifoOut[0][13];
              muxOutConnector[16] = fifoOut[1][13];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[34][9];
              muxOutConnector[27] = fifoOut[35][9];
              muxOutConnector[28] = fifoOut[36][9];
              muxOutConnector[29] = fifoOut[37][9];
              muxOutConnector[30] = fifoOut[38][9];
              muxOutConnector[31] = fifoOut[39][9];
              muxOutConnector[32] = fifoOut[40][9];
              muxOutConnector[33] = fifoOut[41][9];
              muxOutConnector[34] = fifoOut[42][9];
              muxOutConnector[35] = fifoOut[43][9];
              muxOutConnector[36] = fifoOut[44][9];
              muxOutConnector[37] = fifoOut[45][9];
              muxOutConnector[38] = fifoOut[46][9];
              muxOutConnector[39] = fifoOut[47][9];
              muxOutConnector[40] = fifoOut[48][9];
              muxOutConnector[41] = fifoOut[49][9];
              muxOutConnector[42] = fifoOut[50][9];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
