`timescale 1ns / 1ps
module LMem0To1_511_circ9_ys_scripted(
        muxOut,
        ly0In,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 11;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

reg   feedback_en;
reg [ w - 1 : 0 ]column_1[ r - 1 : 0 ];
reg chip_en;
wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(chip_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= column_1[i];
         end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
  feedback_en=rd_en;
      if(wr_en)begin
        chip_en=wr_en;
      end
      else begin
        chip_en=feedback_en;
      end
   if(feedback_en)begin
      for(i = r-1; i > -1; i=i-1) begin
        column_1[i] <= fifoOut[i][c-1];
      end
   end
   else begin
      for(i = r-1; i > -1; i=i-1) begin
        column_1[i] <= ly0InConnector[i];
      end
    end
end
always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[15][10];
              muxOutConnector[1] = fifoOut[16][10];
              muxOutConnector[2] = fifoOut[17][10];
              muxOutConnector[3] = fifoOut[18][10];
              muxOutConnector[4] = fifoOut[19][10];
              muxOutConnector[5] = fifoOut[20][10];
              muxOutConnector[6] = fifoOut[21][10];
              muxOutConnector[7] = fifoOut[22][10];
              muxOutConnector[8] = fifoOut[23][10];
              muxOutConnector[9] = fifoOut[24][10];
              muxOutConnector[10] = fifoOut[25][10];
              muxOutConnector[11] = fifoOut[0][9];
              muxOutConnector[12] = fifoOut[1][9];
              muxOutConnector[13] = fifoOut[2][9];
              muxOutConnector[14] = fifoOut[3][9];
              muxOutConnector[15] = fifoOut[4][9];
              muxOutConnector[16] = fifoOut[5][9];
              muxOutConnector[17] = fifoOut[6][9];
              muxOutConnector[18] = fifoOut[7][9];
              muxOutConnector[19] = fifoOut[8][9];
              muxOutConnector[20] = fifoOut[9][9];
              muxOutConnector[21] = fifoOut[10][9];
              muxOutConnector[22] = fifoOut[11][9];
              muxOutConnector[23] = fifoOut[12][9];
              muxOutConnector[24] = fifoOut[13][9];
              muxOutConnector[25] = fifoOut[14][9];
              muxOutConnector[26] = fifoOut[8][4];
              muxOutConnector[27] = fifoOut[9][4];
              muxOutConnector[28] = fifoOut[10][4];
              muxOutConnector[29] = fifoOut[11][4];
              muxOutConnector[30] = fifoOut[12][4];
              muxOutConnector[31] = fifoOut[13][4];
              muxOutConnector[32] = fifoOut[14][4];
              muxOutConnector[33] = fifoOut[15][4];
              muxOutConnector[34] = fifoOut[16][4];
              muxOutConnector[35] = fifoOut[17][4];
              muxOutConnector[36] = fifoOut[18][4];
              muxOutConnector[37] = fifoOut[19][4];
              muxOutConnector[38] = fifoOut[20][4];
              muxOutConnector[39] = fifoOut[21][4];
              muxOutConnector[40] = fifoOut[22][4];
              muxOutConnector[41] = fifoOut[23][4];
              muxOutConnector[42] = fifoOut[24][4];
              muxOutConnector[43] = fifoOut[25][4];
              muxOutConnector[44] = fifoOut[0][3];
              muxOutConnector[45] = fifoOut[1][3];
              muxOutConnector[46] = fifoOut[2][3];
              muxOutConnector[47] = fifoOut[3][3];
              muxOutConnector[48] = fifoOut[4][3];
              muxOutConnector[49] = fifoOut[5][3];
              muxOutConnector[50] = fifoOut[6][3];
              muxOutConnector[51] = fifoOut[7][3];
       end
       1: begin
              muxOutConnector[0] = fifoOut[15][10];
              muxOutConnector[1] = fifoOut[16][10];
              muxOutConnector[2] = fifoOut[17][10];
              muxOutConnector[3] = fifoOut[18][10];
              muxOutConnector[4] = fifoOut[19][10];
              muxOutConnector[5] = fifoOut[20][10];
              muxOutConnector[6] = fifoOut[21][10];
              muxOutConnector[7] = fifoOut[22][10];
              muxOutConnector[8] = fifoOut[23][10];
              muxOutConnector[9] = fifoOut[24][10];
              muxOutConnector[10] = fifoOut[25][10];
              muxOutConnector[11] = fifoOut[0][9];
              muxOutConnector[12] = fifoOut[1][9];
              muxOutConnector[13] = fifoOut[2][9];
              muxOutConnector[14] = fifoOut[3][9];
              muxOutConnector[15] = fifoOut[4][9];
              muxOutConnector[16] = fifoOut[5][9];
              muxOutConnector[17] = fifoOut[6][9];
              muxOutConnector[18] = fifoOut[7][9];
              muxOutConnector[19] = fifoOut[8][9];
              muxOutConnector[20] = fifoOut[9][9];
              muxOutConnector[21] = fifoOut[10][9];
              muxOutConnector[22] = fifoOut[11][9];
              muxOutConnector[23] = fifoOut[12][9];
              muxOutConnector[24] = fifoOut[13][9];
              muxOutConnector[25] = fifoOut[14][9];
              muxOutConnector[26] = fifoOut[8][4];
              muxOutConnector[27] = fifoOut[9][4];
              muxOutConnector[28] = fifoOut[10][4];
              muxOutConnector[29] = fifoOut[11][4];
              muxOutConnector[30] = fifoOut[12][4];
              muxOutConnector[31] = fifoOut[13][4];
              muxOutConnector[32] = fifoOut[14][4];
              muxOutConnector[33] = fifoOut[15][4];
              muxOutConnector[34] = fifoOut[16][4];
              muxOutConnector[35] = fifoOut[17][4];
              muxOutConnector[36] = fifoOut[18][4];
              muxOutConnector[37] = fifoOut[19][4];
              muxOutConnector[38] = fifoOut[20][4];
              muxOutConnector[39] = fifoOut[21][4];
              muxOutConnector[40] = fifoOut[22][4];
              muxOutConnector[41] = fifoOut[23][4];
              muxOutConnector[42] = fifoOut[24][4];
              muxOutConnector[43] = fifoOut[25][4];
              muxOutConnector[44] = fifoOut[0][3];
              muxOutConnector[45] = fifoOut[1][3];
              muxOutConnector[46] = fifoOut[2][3];
              muxOutConnector[47] = fifoOut[3][3];
              muxOutConnector[48] = fifoOut[4][3];
              muxOutConnector[49] = fifoOut[5][3];
              muxOutConnector[50] = fifoOut[6][3];
              muxOutConnector[51] = fifoOut[7][3];
       end
       2: begin
              muxOutConnector[0] = fifoOut[15][10];
              muxOutConnector[1] = fifoOut[16][10];
              muxOutConnector[2] = fifoOut[17][10];
              muxOutConnector[3] = fifoOut[18][10];
              muxOutConnector[4] = fifoOut[19][10];
              muxOutConnector[5] = fifoOut[20][10];
              muxOutConnector[6] = fifoOut[21][10];
              muxOutConnector[7] = fifoOut[22][10];
              muxOutConnector[8] = fifoOut[23][10];
              muxOutConnector[9] = fifoOut[24][10];
              muxOutConnector[10] = fifoOut[25][10];
              muxOutConnector[11] = fifoOut[0][9];
              muxOutConnector[12] = fifoOut[1][9];
              muxOutConnector[13] = fifoOut[2][9];
              muxOutConnector[14] = fifoOut[3][9];
              muxOutConnector[15] = fifoOut[4][9];
              muxOutConnector[16] = fifoOut[5][9];
              muxOutConnector[17] = fifoOut[6][9];
              muxOutConnector[18] = fifoOut[7][9];
              muxOutConnector[19] = fifoOut[8][9];
              muxOutConnector[20] = fifoOut[9][9];
              muxOutConnector[21] = fifoOut[10][9];
              muxOutConnector[22] = fifoOut[11][9];
              muxOutConnector[23] = fifoOut[12][9];
              muxOutConnector[24] = fifoOut[13][9];
              muxOutConnector[25] = fifoOut[14][9];
              muxOutConnector[26] = fifoOut[8][4];
              muxOutConnector[27] = fifoOut[9][4];
              muxOutConnector[28] = fifoOut[10][4];
              muxOutConnector[29] = fifoOut[11][4];
              muxOutConnector[30] = fifoOut[12][4];
              muxOutConnector[31] = fifoOut[13][4];
              muxOutConnector[32] = fifoOut[14][4];
              muxOutConnector[33] = fifoOut[15][4];
              muxOutConnector[34] = fifoOut[16][4];
              muxOutConnector[35] = fifoOut[17][4];
              muxOutConnector[36] = fifoOut[18][4];
              muxOutConnector[37] = fifoOut[19][4];
              muxOutConnector[38] = fifoOut[20][4];
              muxOutConnector[39] = fifoOut[21][4];
              muxOutConnector[40] = fifoOut[22][4];
              muxOutConnector[41] = fifoOut[23][4];
              muxOutConnector[42] = fifoOut[24][4];
              muxOutConnector[43] = fifoOut[25][4];
              muxOutConnector[44] = fifoOut[0][3];
              muxOutConnector[45] = fifoOut[1][3];
              muxOutConnector[46] = fifoOut[2][3];
              muxOutConnector[47] = fifoOut[3][3];
              muxOutConnector[48] = fifoOut[4][3];
              muxOutConnector[49] = fifoOut[5][3];
              muxOutConnector[50] = fifoOut[6][3];
              muxOutConnector[51] = fifoOut[7][3];
       end
       3: begin
              muxOutConnector[0] = fifoOut[15][10];
              muxOutConnector[1] = fifoOut[16][10];
              muxOutConnector[2] = fifoOut[17][10];
              muxOutConnector[3] = fifoOut[18][10];
              muxOutConnector[4] = fifoOut[19][10];
              muxOutConnector[5] = fifoOut[20][10];
              muxOutConnector[6] = fifoOut[21][10];
              muxOutConnector[7] = fifoOut[22][10];
              muxOutConnector[8] = fifoOut[23][10];
              muxOutConnector[9] = fifoOut[24][10];
              muxOutConnector[10] = fifoOut[25][10];
              muxOutConnector[11] = fifoOut[0][9];
              muxOutConnector[12] = fifoOut[1][9];
              muxOutConnector[13] = fifoOut[2][9];
              muxOutConnector[14] = fifoOut[3][9];
              muxOutConnector[15] = fifoOut[4][9];
              muxOutConnector[16] = fifoOut[5][9];
              muxOutConnector[17] = fifoOut[6][9];
              muxOutConnector[18] = fifoOut[7][9];
              muxOutConnector[19] = fifoOut[8][9];
              muxOutConnector[20] = fifoOut[9][9];
              muxOutConnector[21] = fifoOut[10][9];
              muxOutConnector[22] = fifoOut[11][9];
              muxOutConnector[23] = fifoOut[12][9];
              muxOutConnector[24] = fifoOut[13][9];
              muxOutConnector[25] = fifoOut[14][9];
              muxOutConnector[26] = fifoOut[8][4];
              muxOutConnector[27] = fifoOut[9][4];
              muxOutConnector[28] = fifoOut[10][4];
              muxOutConnector[29] = fifoOut[11][4];
              muxOutConnector[30] = fifoOut[12][4];
              muxOutConnector[31] = fifoOut[13][4];
              muxOutConnector[32] = fifoOut[14][4];
              muxOutConnector[33] = fifoOut[15][4];
              muxOutConnector[34] = fifoOut[16][4];
              muxOutConnector[35] = fifoOut[17][4];
              muxOutConnector[36] = fifoOut[18][4];
              muxOutConnector[37] = fifoOut[19][4];
              muxOutConnector[38] = fifoOut[20][4];
              muxOutConnector[39] = fifoOut[21][4];
              muxOutConnector[40] = fifoOut[22][4];
              muxOutConnector[41] = fifoOut[23][4];
              muxOutConnector[42] = fifoOut[24][4];
              muxOutConnector[43] = fifoOut[25][4];
              muxOutConnector[44] = fifoOut[0][3];
              muxOutConnector[45] = fifoOut[1][3];
              muxOutConnector[46] = fifoOut[2][3];
              muxOutConnector[47] = fifoOut[3][3];
              muxOutConnector[48] = fifoOut[4][3];
              muxOutConnector[49] = fifoOut[5][3];
              muxOutConnector[50] = fifoOut[6][3];
              muxOutConnector[51] = fifoOut[7][3];
       end
       4: begin
              muxOutConnector[0] = fifoOut[15][10];
              muxOutConnector[1] = fifoOut[16][10];
              muxOutConnector[2] = fifoOut[17][10];
              muxOutConnector[3] = fifoOut[18][10];
              muxOutConnector[4] = fifoOut[19][10];
              muxOutConnector[5] = fifoOut[20][10];
              muxOutConnector[6] = fifoOut[21][10];
              muxOutConnector[7] = fifoOut[22][10];
              muxOutConnector[8] = fifoOut[23][10];
              muxOutConnector[9] = fifoOut[24][10];
              muxOutConnector[10] = fifoOut[25][10];
              muxOutConnector[11] = fifoOut[0][9];
              muxOutConnector[12] = fifoOut[1][9];
              muxOutConnector[13] = fifoOut[2][9];
              muxOutConnector[14] = fifoOut[3][9];
              muxOutConnector[15] = fifoOut[4][9];
              muxOutConnector[16] = fifoOut[5][9];
              muxOutConnector[17] = fifoOut[6][9];
              muxOutConnector[18] = fifoOut[7][9];
              muxOutConnector[19] = fifoOut[8][9];
              muxOutConnector[20] = fifoOut[9][9];
              muxOutConnector[21] = fifoOut[10][9];
              muxOutConnector[22] = fifoOut[11][9];
              muxOutConnector[23] = fifoOut[12][9];
              muxOutConnector[24] = fifoOut[13][9];
              muxOutConnector[25] = fifoOut[14][9];
              muxOutConnector[26] = fifoOut[8][4];
              muxOutConnector[27] = fifoOut[9][4];
              muxOutConnector[28] = fifoOut[10][4];
              muxOutConnector[29] = fifoOut[11][4];
              muxOutConnector[30] = fifoOut[12][4];
              muxOutConnector[31] = fifoOut[13][4];
              muxOutConnector[32] = fifoOut[14][4];
              muxOutConnector[33] = fifoOut[15][4];
              muxOutConnector[34] = fifoOut[16][4];
              muxOutConnector[35] = fifoOut[27][3];
              muxOutConnector[36] = fifoOut[28][3];
              muxOutConnector[37] = fifoOut[29][3];
              muxOutConnector[38] = fifoOut[30][3];
              muxOutConnector[39] = fifoOut[31][3];
              muxOutConnector[40] = fifoOut[32][3];
              muxOutConnector[41] = fifoOut[33][3];
              muxOutConnector[42] = fifoOut[34][3];
              muxOutConnector[43] = fifoOut[35][3];
              muxOutConnector[44] = fifoOut[36][3];
              muxOutConnector[45] = fifoOut[37][3];
              muxOutConnector[46] = fifoOut[38][3];
              muxOutConnector[47] = fifoOut[39][3];
              muxOutConnector[48] = fifoOut[40][3];
              muxOutConnector[49] = fifoOut[41][3];
              muxOutConnector[50] = fifoOut[42][3];
              muxOutConnector[51] = fifoOut[43][3];
       end
       5: begin
              muxOutConnector[0] = fifoOut[15][10];
              muxOutConnector[1] = fifoOut[16][10];
              muxOutConnector[2] = fifoOut[17][10];
              muxOutConnector[3] = fifoOut[18][10];
              muxOutConnector[4] = fifoOut[19][10];
              muxOutConnector[5] = fifoOut[20][10];
              muxOutConnector[6] = fifoOut[21][10];
              muxOutConnector[7] = fifoOut[22][10];
              muxOutConnector[8] = fifoOut[23][10];
              muxOutConnector[9] = fifoOut[24][10];
              muxOutConnector[10] = fifoOut[25][10];
              muxOutConnector[11] = fifoOut[0][9];
              muxOutConnector[12] = fifoOut[1][9];
              muxOutConnector[13] = fifoOut[2][9];
              muxOutConnector[14] = fifoOut[3][9];
              muxOutConnector[15] = fifoOut[4][9];
              muxOutConnector[16] = fifoOut[5][9];
              muxOutConnector[17] = fifoOut[6][9];
              muxOutConnector[18] = fifoOut[7][9];
              muxOutConnector[19] = fifoOut[8][9];
              muxOutConnector[20] = fifoOut[9][9];
              muxOutConnector[21] = fifoOut[10][9];
              muxOutConnector[22] = fifoOut[11][9];
              muxOutConnector[23] = fifoOut[12][9];
              muxOutConnector[24] = fifoOut[13][9];
              muxOutConnector[25] = fifoOut[14][9];
              muxOutConnector[26] = fifoOut[44][4];
              muxOutConnector[27] = fifoOut[45][4];
              muxOutConnector[28] = fifoOut[46][4];
              muxOutConnector[29] = fifoOut[47][4];
              muxOutConnector[30] = fifoOut[48][4];
              muxOutConnector[31] = fifoOut[49][4];
              muxOutConnector[32] = fifoOut[50][4];
              muxOutConnector[33] = fifoOut[51][4];
              muxOutConnector[34] = fifoOut[26][3];
              muxOutConnector[35] = fifoOut[27][3];
              muxOutConnector[36] = fifoOut[28][3];
              muxOutConnector[37] = fifoOut[29][3];
              muxOutConnector[38] = fifoOut[30][3];
              muxOutConnector[39] = fifoOut[31][3];
              muxOutConnector[40] = fifoOut[32][3];
              muxOutConnector[41] = fifoOut[33][3];
              muxOutConnector[42] = fifoOut[34][3];
              muxOutConnector[43] = fifoOut[35][3];
              muxOutConnector[44] = fifoOut[36][3];
              muxOutConnector[45] = fifoOut[37][3];
              muxOutConnector[46] = fifoOut[38][3];
              muxOutConnector[47] = fifoOut[39][3];
              muxOutConnector[48] = fifoOut[40][3];
              muxOutConnector[49] = fifoOut[41][3];
              muxOutConnector[50] = fifoOut[42][3];
              muxOutConnector[51] = fifoOut[43][3];
       end
       6: begin
              muxOutConnector[0] = fifoOut[15][10];
              muxOutConnector[1] = fifoOut[16][10];
              muxOutConnector[2] = fifoOut[17][10];
              muxOutConnector[3] = fifoOut[18][10];
              muxOutConnector[4] = fifoOut[19][10];
              muxOutConnector[5] = fifoOut[20][10];
              muxOutConnector[6] = fifoOut[21][10];
              muxOutConnector[7] = fifoOut[22][10];
              muxOutConnector[8] = fifoOut[23][10];
              muxOutConnector[9] = fifoOut[24][10];
              muxOutConnector[10] = fifoOut[25][10];
              muxOutConnector[11] = fifoOut[0][9];
              muxOutConnector[12] = fifoOut[1][9];
              muxOutConnector[13] = fifoOut[2][9];
              muxOutConnector[14] = fifoOut[3][9];
              muxOutConnector[15] = fifoOut[4][9];
              muxOutConnector[16] = fifoOut[5][9];
              muxOutConnector[17] = fifoOut[6][9];
              muxOutConnector[18] = fifoOut[7][9];
              muxOutConnector[19] = fifoOut[8][9];
              muxOutConnector[20] = fifoOut[9][9];
              muxOutConnector[21] = fifoOut[10][9];
              muxOutConnector[22] = fifoOut[11][9];
              muxOutConnector[23] = fifoOut[12][9];
              muxOutConnector[24] = fifoOut[13][9];
              muxOutConnector[25] = fifoOut[14][9];
              muxOutConnector[26] = fifoOut[44][4];
              muxOutConnector[27] = fifoOut[45][4];
              muxOutConnector[28] = fifoOut[46][4];
              muxOutConnector[29] = fifoOut[47][4];
              muxOutConnector[30] = fifoOut[48][4];
              muxOutConnector[31] = fifoOut[49][4];
              muxOutConnector[32] = fifoOut[50][4];
              muxOutConnector[33] = fifoOut[51][4];
              muxOutConnector[34] = fifoOut[26][3];
              muxOutConnector[35] = fifoOut[27][3];
              muxOutConnector[36] = fifoOut[28][3];
              muxOutConnector[37] = fifoOut[29][3];
              muxOutConnector[38] = fifoOut[30][3];
              muxOutConnector[39] = fifoOut[31][3];
              muxOutConnector[40] = fifoOut[32][3];
              muxOutConnector[41] = fifoOut[33][3];
              muxOutConnector[42] = fifoOut[34][3];
              muxOutConnector[43] = fifoOut[35][3];
              muxOutConnector[44] = fifoOut[36][3];
              muxOutConnector[45] = fifoOut[37][3];
              muxOutConnector[46] = fifoOut[38][3];
              muxOutConnector[47] = fifoOut[39][3];
              muxOutConnector[48] = fifoOut[40][3];
              muxOutConnector[49] = fifoOut[41][3];
              muxOutConnector[50] = fifoOut[42][3];
              muxOutConnector[51] = fifoOut[43][3];
       end
       7: begin
              muxOutConnector[0] = fifoOut[15][10];
              muxOutConnector[1] = fifoOut[16][10];
              muxOutConnector[2] = fifoOut[17][10];
              muxOutConnector[3] = fifoOut[18][10];
              muxOutConnector[4] = fifoOut[19][10];
              muxOutConnector[5] = fifoOut[20][10];
              muxOutConnector[6] = fifoOut[21][10];
              muxOutConnector[7] = fifoOut[22][10];
              muxOutConnector[8] = fifoOut[23][10];
              muxOutConnector[9] = fifoOut[24][10];
              muxOutConnector[10] = fifoOut[25][10];
              muxOutConnector[11] = fifoOut[0][9];
              muxOutConnector[12] = fifoOut[1][9];
              muxOutConnector[13] = fifoOut[2][9];
              muxOutConnector[14] = fifoOut[3][9];
              muxOutConnector[15] = fifoOut[4][9];
              muxOutConnector[16] = fifoOut[5][9];
              muxOutConnector[17] = fifoOut[6][9];
              muxOutConnector[18] = fifoOut[7][9];
              muxOutConnector[19] = fifoOut[8][9];
              muxOutConnector[20] = fifoOut[9][9];
              muxOutConnector[21] = fifoOut[10][9];
              muxOutConnector[22] = fifoOut[11][9];
              muxOutConnector[23] = fifoOut[12][9];
              muxOutConnector[24] = fifoOut[13][9];
              muxOutConnector[25] = fifoOut[14][9];
              muxOutConnector[26] = fifoOut[44][4];
              muxOutConnector[27] = fifoOut[45][4];
              muxOutConnector[28] = fifoOut[46][4];
              muxOutConnector[29] = fifoOut[47][4];
              muxOutConnector[30] = fifoOut[48][4];
              muxOutConnector[31] = fifoOut[49][4];
              muxOutConnector[32] = fifoOut[50][4];
              muxOutConnector[33] = fifoOut[51][4];
              muxOutConnector[34] = fifoOut[26][3];
              muxOutConnector[35] = fifoOut[27][3];
              muxOutConnector[36] = fifoOut[28][3];
              muxOutConnector[37] = fifoOut[29][3];
              muxOutConnector[38] = fifoOut[30][3];
              muxOutConnector[39] = fifoOut[31][3];
              muxOutConnector[40] = fifoOut[32][3];
              muxOutConnector[41] = fifoOut[33][3];
              muxOutConnector[42] = fifoOut[34][3];
              muxOutConnector[43] = fifoOut[35][3];
              muxOutConnector[44] = fifoOut[36][3];
              muxOutConnector[45] = fifoOut[37][3];
              muxOutConnector[46] = fifoOut[38][3];
              muxOutConnector[47] = fifoOut[39][3];
              muxOutConnector[48] = fifoOut[40][3];
              muxOutConnector[49] = fifoOut[41][3];
              muxOutConnector[50] = fifoOut[42][3];
              muxOutConnector[51] = fifoOut[43][3];
       end
       8: begin
              muxOutConnector[0] = fifoOut[15][10];
              muxOutConnector[1] = fifoOut[16][10];
              muxOutConnector[2] = fifoOut[17][10];
              muxOutConnector[3] = fifoOut[18][10];
              muxOutConnector[4] = fifoOut[19][10];
              muxOutConnector[5] = fifoOut[20][10];
              muxOutConnector[6] = fifoOut[21][10];
              muxOutConnector[7] = fifoOut[22][10];
              muxOutConnector[8] = fifoOut[23][10];
              muxOutConnector[9] = fifoOut[24][10];
              muxOutConnector[10] = fifoOut[25][10];
              muxOutConnector[11] = fifoOut[0][9];
              muxOutConnector[12] = fifoOut[1][9];
              muxOutConnector[13] = fifoOut[2][9];
              muxOutConnector[14] = fifoOut[3][9];
              muxOutConnector[15] = fifoOut[4][9];
              muxOutConnector[16] = fifoOut[5][9];
              muxOutConnector[17] = fifoOut[6][9];
              muxOutConnector[18] = fifoOut[7][9];
              muxOutConnector[19] = fifoOut[8][9];
              muxOutConnector[20] = fifoOut[9][9];
              muxOutConnector[21] = fifoOut[10][9];
              muxOutConnector[22] = fifoOut[11][9];
              muxOutConnector[23] = fifoOut[12][9];
              muxOutConnector[24] = fifoOut[13][9];
              muxOutConnector[25] = fifoOut[14][9];
              muxOutConnector[26] = fifoOut[44][4];
              muxOutConnector[27] = fifoOut[45][4];
              muxOutConnector[28] = fifoOut[46][4];
              muxOutConnector[29] = fifoOut[47][4];
              muxOutConnector[30] = fifoOut[48][4];
              muxOutConnector[31] = fifoOut[49][4];
              muxOutConnector[32] = fifoOut[50][4];
              muxOutConnector[33] = fifoOut[51][4];
              muxOutConnector[34] = fifoOut[26][3];
              muxOutConnector[35] = fifoOut[27][3];
              muxOutConnector[36] = fifoOut[28][3];
              muxOutConnector[37] = fifoOut[29][3];
              muxOutConnector[38] = fifoOut[30][3];
              muxOutConnector[39] = fifoOut[31][3];
              muxOutConnector[40] = fifoOut[32][3];
              muxOutConnector[41] = fifoOut[33][3];
              muxOutConnector[42] = fifoOut[34][3];
              muxOutConnector[43] = fifoOut[35][3];
              muxOutConnector[44] = fifoOut[36][3];
              muxOutConnector[45] = fifoOut[37][3];
              muxOutConnector[46] = fifoOut[38][3];
              muxOutConnector[47] = fifoOut[39][3];
              muxOutConnector[48] = fifoOut[40][3];
              muxOutConnector[49] = fifoOut[41][3];
              muxOutConnector[50] = fifoOut[42][3];
              muxOutConnector[51] = fifoOut[43][3];
       end
       9: begin
              muxOutConnector[0] = fifoOut[15][10];
              muxOutConnector[1] = fifoOut[16][10];
              muxOutConnector[2] = fifoOut[17][10];
              muxOutConnector[3] = fifoOut[18][10];
              muxOutConnector[4] = fifoOut[19][10];
              muxOutConnector[5] = fifoOut[20][10];
              muxOutConnector[6] = fifoOut[21][10];
              muxOutConnector[7] = fifoOut[22][10];
              muxOutConnector[8] = fifoOut[23][10];
              muxOutConnector[9] = fifoOut[24][10];
              muxOutConnector[10] = fifoOut[25][10];
              muxOutConnector[11] = fifoOut[0][9];
              muxOutConnector[12] = fifoOut[1][9];
              muxOutConnector[13] = fifoOut[2][9];
              muxOutConnector[14] = fifoOut[3][9];
              muxOutConnector[15] = fifoOut[4][9];
              muxOutConnector[16] = fifoOut[5][9];
              muxOutConnector[17] = fifoOut[6][9];
              muxOutConnector[18] = fifoOut[7][9];
              muxOutConnector[19] = fifoOut[8][9];
              muxOutConnector[20] = fifoOut[9][9];
              muxOutConnector[21] = fifoOut[10][9];
              muxOutConnector[22] = fifoOut[11][9];
              muxOutConnector[23] = fifoOut[12][9];
              muxOutConnector[24] = fifoOut[13][9];
              muxOutConnector[25] = fifoOut[14][9];
              muxOutConnector[26] = fifoOut[44][4];
              muxOutConnector[27] = fifoOut[45][4];
              muxOutConnector[28] = fifoOut[46][4];
              muxOutConnector[29] = fifoOut[47][4];
              muxOutConnector[30] = fifoOut[48][4];
              muxOutConnector[31] = fifoOut[49][4];
              muxOutConnector[32] = fifoOut[50][4];
              muxOutConnector[33] = fifoOut[51][4];
              muxOutConnector[34] = fifoOut[26][3];
              muxOutConnector[35] = fifoOut[27][3];
              muxOutConnector[36] = fifoOut[28][3];
              muxOutConnector[37] = fifoOut[29][3];
              muxOutConnector[38] = fifoOut[30][3];
              muxOutConnector[39] = fifoOut[31][3];
              muxOutConnector[40] = fifoOut[32][3];
              muxOutConnector[41] = fifoOut[33][3];
              muxOutConnector[42] = fifoOut[34][3];
              muxOutConnector[43] = fifoOut[35][3];
              muxOutConnector[44] = fifoOut[36][3];
              muxOutConnector[45] = fifoOut[37][3];
              muxOutConnector[46] = fifoOut[38][3];
              muxOutConnector[47] = fifoOut[39][3];
              muxOutConnector[48] = fifoOut[40][3];
              muxOutConnector[49] = fifoOut[41][3];
              muxOutConnector[50] = fifoOut[42][3];
              muxOutConnector[51] = fifoOut[43][3];
       end
       10: begin
              muxOutConnector[0] = fifoOut[15][10];
              muxOutConnector[1] = fifoOut[16][10];
              muxOutConnector[2] = fifoOut[27][9];
              muxOutConnector[3] = fifoOut[28][9];
              muxOutConnector[4] = fifoOut[29][9];
              muxOutConnector[5] = fifoOut[30][9];
              muxOutConnector[6] = fifoOut[31][9];
              muxOutConnector[7] = fifoOut[32][9];
              muxOutConnector[8] = fifoOut[33][9];
              muxOutConnector[9] = fifoOut[34][9];
              muxOutConnector[10] = fifoOut[35][9];
              muxOutConnector[11] = fifoOut[36][9];
              muxOutConnector[12] = fifoOut[37][9];
              muxOutConnector[13] = fifoOut[38][9];
              muxOutConnector[14] = fifoOut[39][9];
              muxOutConnector[15] = fifoOut[40][9];
              muxOutConnector[16] = fifoOut[41][9];
              muxOutConnector[17] = fifoOut[42][9];
              muxOutConnector[18] = fifoOut[43][9];
              muxOutConnector[19] = fifoOut[44][9];
              muxOutConnector[20] = fifoOut[45][9];
              muxOutConnector[21] = fifoOut[46][9];
              muxOutConnector[22] = fifoOut[47][9];
              muxOutConnector[23] = fifoOut[48][9];
              muxOutConnector[24] = fifoOut[49][9];
              muxOutConnector[25] = fifoOut[50][9];
              muxOutConnector[26] = fifoOut[44][4];
              muxOutConnector[27] = fifoOut[45][4];
              muxOutConnector[28] = fifoOut[46][4];
              muxOutConnector[29] = fifoOut[47][4];
              muxOutConnector[30] = fifoOut[48][4];
              muxOutConnector[31] = fifoOut[49][4];
              muxOutConnector[32] = fifoOut[50][4];
              muxOutConnector[33] = fifoOut[51][4];
              muxOutConnector[34] = fifoOut[26][3];
              muxOutConnector[35] = fifoOut[27][3];
              muxOutConnector[36] = fifoOut[28][3];
              muxOutConnector[37] = fifoOut[29][3];
              muxOutConnector[38] = fifoOut[30][3];
              muxOutConnector[39] = fifoOut[31][3];
              muxOutConnector[40] = fifoOut[32][3];
              muxOutConnector[41] = fifoOut[33][3];
              muxOutConnector[42] = fifoOut[34][3];
              muxOutConnector[43] = fifoOut[35][3];
              muxOutConnector[44] = fifoOut[36][3];
              muxOutConnector[45] = fifoOut[37][3];
              muxOutConnector[46] = fifoOut[38][3];
              muxOutConnector[47] = fifoOut[39][3];
              muxOutConnector[48] = fifoOut[40][3];
              muxOutConnector[49] = fifoOut[41][3];
              muxOutConnector[50] = fifoOut[42][3];
              muxOutConnector[51] = fifoOut[43][3];
       end
       11: begin
              muxOutConnector[0] = fifoOut[51][10];
              muxOutConnector[1] = fifoOut[26][9];
              muxOutConnector[2] = fifoOut[27][9];
              muxOutConnector[3] = fifoOut[28][9];
              muxOutConnector[4] = fifoOut[29][9];
              muxOutConnector[5] = fifoOut[30][9];
              muxOutConnector[6] = fifoOut[31][9];
              muxOutConnector[7] = fifoOut[32][9];
              muxOutConnector[8] = fifoOut[33][9];
              muxOutConnector[9] = fifoOut[34][9];
              muxOutConnector[10] = fifoOut[35][9];
              muxOutConnector[11] = fifoOut[36][9];
              muxOutConnector[12] = fifoOut[37][9];
              muxOutConnector[13] = fifoOut[38][9];
              muxOutConnector[14] = fifoOut[39][9];
              muxOutConnector[15] = fifoOut[40][9];
              muxOutConnector[16] = fifoOut[41][9];
              muxOutConnector[17] = fifoOut[42][9];
              muxOutConnector[18] = fifoOut[43][9];
              muxOutConnector[19] = fifoOut[44][9];
              muxOutConnector[20] = fifoOut[45][9];
              muxOutConnector[21] = fifoOut[46][9];
              muxOutConnector[22] = fifoOut[47][9];
              muxOutConnector[23] = fifoOut[48][9];
              muxOutConnector[24] = fifoOut[49][9];
              muxOutConnector[25] = fifoOut[50][9];
              muxOutConnector[26] = fifoOut[44][4];
              muxOutConnector[27] = fifoOut[45][4];
              muxOutConnector[28] = fifoOut[46][4];
              muxOutConnector[29] = fifoOut[47][4];
              muxOutConnector[30] = fifoOut[48][4];
              muxOutConnector[31] = fifoOut[49][4];
              muxOutConnector[32] = fifoOut[50][4];
              muxOutConnector[33] = fifoOut[51][4];
              muxOutConnector[34] = fifoOut[26][3];
              muxOutConnector[35] = fifoOut[27][3];
              muxOutConnector[36] = fifoOut[28][3];
              muxOutConnector[37] = fifoOut[29][3];
              muxOutConnector[38] = fifoOut[30][3];
              muxOutConnector[39] = fifoOut[31][3];
              muxOutConnector[40] = fifoOut[32][3];
              muxOutConnector[41] = fifoOut[33][3];
              muxOutConnector[42] = fifoOut[34][3];
              muxOutConnector[43] = fifoOut[35][3];
              muxOutConnector[44] = fifoOut[36][3];
              muxOutConnector[45] = fifoOut[37][3];
              muxOutConnector[46] = fifoOut[38][3];
              muxOutConnector[47] = fifoOut[39][3];
              muxOutConnector[48] = fifoOut[40][3];
              muxOutConnector[49] = fifoOut[41][3];
              muxOutConnector[50] = fifoOut[42][3];
              muxOutConnector[51] = fifoOut[43][3];
       end
       12: begin
              muxOutConnector[0] = fifoOut[51][10];
              muxOutConnector[1] = fifoOut[26][9];
              muxOutConnector[2] = fifoOut[27][9];
              muxOutConnector[3] = fifoOut[28][9];
              muxOutConnector[4] = fifoOut[29][9];
              muxOutConnector[5] = fifoOut[30][9];
              muxOutConnector[6] = fifoOut[31][9];
              muxOutConnector[7] = fifoOut[32][9];
              muxOutConnector[8] = fifoOut[33][9];
              muxOutConnector[9] = fifoOut[34][9];
              muxOutConnector[10] = fifoOut[35][9];
              muxOutConnector[11] = fifoOut[36][9];
              muxOutConnector[12] = fifoOut[37][9];
              muxOutConnector[13] = fifoOut[38][9];
              muxOutConnector[14] = fifoOut[39][9];
              muxOutConnector[15] = fifoOut[40][9];
              muxOutConnector[16] = fifoOut[41][9];
              muxOutConnector[17] = fifoOut[42][9];
              muxOutConnector[18] = fifoOut[43][9];
              muxOutConnector[19] = fifoOut[44][9];
              muxOutConnector[20] = fifoOut[45][9];
              muxOutConnector[21] = fifoOut[46][9];
              muxOutConnector[22] = fifoOut[47][9];
              muxOutConnector[23] = fifoOut[48][9];
              muxOutConnector[24] = fifoOut[49][9];
              muxOutConnector[25] = fifoOut[50][9];
              muxOutConnector[26] = fifoOut[44][4];
              muxOutConnector[27] = fifoOut[45][4];
              muxOutConnector[28] = fifoOut[46][4];
              muxOutConnector[29] = fifoOut[47][4];
              muxOutConnector[30] = fifoOut[48][4];
              muxOutConnector[31] = fifoOut[49][4];
              muxOutConnector[32] = fifoOut[50][4];
              muxOutConnector[33] = fifoOut[51][4];
              muxOutConnector[34] = fifoOut[26][3];
              muxOutConnector[35] = fifoOut[27][3];
              muxOutConnector[36] = fifoOut[28][3];
              muxOutConnector[37] = fifoOut[29][3];
              muxOutConnector[38] = fifoOut[30][3];
              muxOutConnector[39] = fifoOut[31][3];
              muxOutConnector[40] = fifoOut[32][3];
              muxOutConnector[41] = fifoOut[33][3];
              muxOutConnector[42] = fifoOut[34][3];
              muxOutConnector[43] = fifoOut[35][3];
              muxOutConnector[44] = fifoOut[36][3];
              muxOutConnector[45] = fifoOut[37][3];
              muxOutConnector[46] = fifoOut[38][3];
              muxOutConnector[47] = fifoOut[39][3];
              muxOutConnector[48] = fifoOut[40][3];
              muxOutConnector[49] = fifoOut[41][3];
              muxOutConnector[50] = fifoOut[42][3];
              muxOutConnector[51] = fifoOut[43][3];
       end
       13: begin
              muxOutConnector[0] = fifoOut[51][10];
              muxOutConnector[1] = fifoOut[26][9];
              muxOutConnector[2] = fifoOut[27][9];
              muxOutConnector[3] = fifoOut[28][9];
              muxOutConnector[4] = fifoOut[29][9];
              muxOutConnector[5] = fifoOut[30][9];
              muxOutConnector[6] = fifoOut[31][9];
              muxOutConnector[7] = fifoOut[32][9];
              muxOutConnector[8] = fifoOut[33][9];
              muxOutConnector[9] = fifoOut[34][9];
              muxOutConnector[10] = fifoOut[35][9];
              muxOutConnector[11] = fifoOut[36][9];
              muxOutConnector[12] = fifoOut[37][9];
              muxOutConnector[13] = fifoOut[38][9];
              muxOutConnector[14] = fifoOut[39][9];
              muxOutConnector[15] = fifoOut[40][9];
              muxOutConnector[16] = fifoOut[41][9];
              muxOutConnector[17] = fifoOut[42][9];
              muxOutConnector[18] = fifoOut[43][9];
              muxOutConnector[19] = fifoOut[44][9];
              muxOutConnector[20] = fifoOut[45][9];
              muxOutConnector[21] = fifoOut[46][9];
              muxOutConnector[22] = fifoOut[47][9];
              muxOutConnector[23] = fifoOut[48][9];
              muxOutConnector[24] = fifoOut[49][9];
              muxOutConnector[25] = fifoOut[50][9];
              muxOutConnector[26] = fifoOut[44][4];
              muxOutConnector[27] = fifoOut[45][4];
              muxOutConnector[28] = fifoOut[46][4];
              muxOutConnector[29] = fifoOut[47][4];
              muxOutConnector[30] = fifoOut[48][4];
              muxOutConnector[31] = fifoOut[49][4];
              muxOutConnector[32] = fifoOut[50][4];
              muxOutConnector[33] = fifoOut[51][4];
              muxOutConnector[34] = fifoOut[26][3];
              muxOutConnector[35] = fifoOut[27][3];
              muxOutConnector[36] = fifoOut[28][3];
              muxOutConnector[37] = fifoOut[29][3];
              muxOutConnector[38] = fifoOut[30][3];
              muxOutConnector[39] = fifoOut[31][3];
              muxOutConnector[40] = fifoOut[32][3];
              muxOutConnector[41] = fifoOut[33][3];
              muxOutConnector[42] = fifoOut[34][3];
              muxOutConnector[43] = fifoOut[35][3];
              muxOutConnector[44] = fifoOut[36][3];
              muxOutConnector[45] = fifoOut[37][3];
              muxOutConnector[46] = fifoOut[38][3];
              muxOutConnector[47] = fifoOut[39][3];
              muxOutConnector[48] = fifoOut[40][3];
              muxOutConnector[49] = fifoOut[41][3];
              muxOutConnector[50] = fifoOut[42][3];
              muxOutConnector[51] = fifoOut[43][3];
       end
       14: begin
              muxOutConnector[0] = fifoOut[51][10];
              muxOutConnector[1] = fifoOut[26][9];
              muxOutConnector[2] = fifoOut[27][9];
              muxOutConnector[3] = fifoOut[28][9];
              muxOutConnector[4] = fifoOut[29][9];
              muxOutConnector[5] = fifoOut[30][9];
              muxOutConnector[6] = fifoOut[31][9];
              muxOutConnector[7] = fifoOut[32][9];
              muxOutConnector[8] = fifoOut[33][9];
              muxOutConnector[9] = fifoOut[34][9];
              muxOutConnector[10] = fifoOut[35][9];
              muxOutConnector[11] = fifoOut[36][9];
              muxOutConnector[12] = fifoOut[37][9];
              muxOutConnector[13] = fifoOut[38][9];
              muxOutConnector[14] = fifoOut[39][9];
              muxOutConnector[15] = fifoOut[40][9];
              muxOutConnector[16] = fifoOut[41][9];
              muxOutConnector[17] = fifoOut[42][9];
              muxOutConnector[18] = fifoOut[43][9];
              muxOutConnector[19] = fifoOut[44][9];
              muxOutConnector[20] = fifoOut[45][9];
              muxOutConnector[21] = fifoOut[46][9];
              muxOutConnector[22] = fifoOut[47][9];
              muxOutConnector[23] = fifoOut[48][9];
              muxOutConnector[24] = fifoOut[49][9];
              muxOutConnector[25] = fifoOut[50][9];
              muxOutConnector[26] = fifoOut[44][4];
              muxOutConnector[27] = fifoOut[45][4];
              muxOutConnector[28] = fifoOut[46][4];
              muxOutConnector[29] = fifoOut[47][4];
              muxOutConnector[30] = fifoOut[48][4];
              muxOutConnector[31] = fifoOut[49][4];
              muxOutConnector[32] = fifoOut[50][4];
              muxOutConnector[33] = fifoOut[51][4];
              muxOutConnector[34] = fifoOut[26][3];
              muxOutConnector[35] = fifoOut[27][3];
              muxOutConnector[36] = fifoOut[28][3];
              muxOutConnector[37] = fifoOut[29][3];
              muxOutConnector[38] = fifoOut[30][3];
              muxOutConnector[39] = fifoOut[31][3];
              muxOutConnector[40] = fifoOut[32][3];
              muxOutConnector[41] = fifoOut[33][3];
              muxOutConnector[42] = fifoOut[34][3];
              muxOutConnector[43] = fifoOut[35][3];
              muxOutConnector[44] = fifoOut[36][3];
              muxOutConnector[45] = fifoOut[37][3];
              muxOutConnector[46] = fifoOut[38][3];
              muxOutConnector[47] = fifoOut[39][3];
              muxOutConnector[48] = fifoOut[40][3];
              muxOutConnector[49] = fifoOut[41][3];
              muxOutConnector[50] = fifoOut[42][3];
              muxOutConnector[51] = fifoOut[16][1];
       end
       15: begin
              muxOutConnector[0] = fifoOut[51][10];
              muxOutConnector[1] = fifoOut[26][9];
              muxOutConnector[2] = fifoOut[27][9];
              muxOutConnector[3] = fifoOut[28][9];
              muxOutConnector[4] = fifoOut[29][9];
              muxOutConnector[5] = fifoOut[30][9];
              muxOutConnector[6] = fifoOut[31][9];
              muxOutConnector[7] = fifoOut[32][9];
              muxOutConnector[8] = fifoOut[33][9];
              muxOutConnector[9] = fifoOut[34][9];
              muxOutConnector[10] = fifoOut[35][9];
              muxOutConnector[11] = fifoOut[36][9];
              muxOutConnector[12] = fifoOut[37][9];
              muxOutConnector[13] = fifoOut[38][9];
              muxOutConnector[14] = fifoOut[39][9];
              muxOutConnector[15] = fifoOut[40][9];
              muxOutConnector[16] = fifoOut[41][9];
              muxOutConnector[17] = fifoOut[42][9];
              muxOutConnector[18] = fifoOut[43][9];
              muxOutConnector[19] = fifoOut[44][9];
              muxOutConnector[20] = fifoOut[45][9];
              muxOutConnector[21] = fifoOut[46][9];
              muxOutConnector[22] = fifoOut[47][9];
              muxOutConnector[23] = fifoOut[48][9];
              muxOutConnector[24] = fifoOut[49][9];
              muxOutConnector[25] = fifoOut[50][9];
              muxOutConnector[26] = fifoOut[17][2];
              muxOutConnector[27] = fifoOut[18][2];
              muxOutConnector[28] = fifoOut[19][2];
              muxOutConnector[29] = fifoOut[20][2];
              muxOutConnector[30] = fifoOut[21][2];
              muxOutConnector[31] = fifoOut[22][2];
              muxOutConnector[32] = fifoOut[23][2];
              muxOutConnector[33] = fifoOut[24][2];
              muxOutConnector[34] = fifoOut[25][2];
              muxOutConnector[35] = fifoOut[0][1];
              muxOutConnector[36] = fifoOut[1][1];
              muxOutConnector[37] = fifoOut[2][1];
              muxOutConnector[38] = fifoOut[3][1];
              muxOutConnector[39] = fifoOut[4][1];
              muxOutConnector[40] = fifoOut[5][1];
              muxOutConnector[41] = fifoOut[6][1];
              muxOutConnector[42] = fifoOut[7][1];
              muxOutConnector[43] = fifoOut[8][1];
              muxOutConnector[44] = fifoOut[9][1];
              muxOutConnector[45] = fifoOut[10][1];
              muxOutConnector[46] = fifoOut[11][1];
              muxOutConnector[47] = fifoOut[12][1];
              muxOutConnector[48] = fifoOut[13][1];
              muxOutConnector[49] = fifoOut[14][1];
              muxOutConnector[50] = fifoOut[15][1];
              muxOutConnector[51] = fifoOut[16][1];
       end
       16: begin
              muxOutConnector[0] = fifoOut[51][10];
              muxOutConnector[1] = fifoOut[26][9];
              muxOutConnector[2] = fifoOut[27][9];
              muxOutConnector[3] = fifoOut[28][9];
              muxOutConnector[4] = fifoOut[29][9];
              muxOutConnector[5] = fifoOut[30][9];
              muxOutConnector[6] = fifoOut[31][9];
              muxOutConnector[7] = fifoOut[32][9];
              muxOutConnector[8] = fifoOut[33][9];
              muxOutConnector[9] = fifoOut[34][9];
              muxOutConnector[10] = fifoOut[35][9];
              muxOutConnector[11] = fifoOut[36][9];
              muxOutConnector[12] = fifoOut[37][9];
              muxOutConnector[13] = fifoOut[38][9];
              muxOutConnector[14] = fifoOut[39][9];
              muxOutConnector[15] = fifoOut[40][9];
              muxOutConnector[16] = fifoOut[41][9];
              muxOutConnector[17] = fifoOut[42][9];
              muxOutConnector[18] = fifoOut[43][9];
              muxOutConnector[19] = fifoOut[44][9];
              muxOutConnector[20] = fifoOut[45][9];
              muxOutConnector[21] = fifoOut[46][9];
              muxOutConnector[22] = fifoOut[47][9];
              muxOutConnector[23] = fifoOut[48][9];
              muxOutConnector[24] = fifoOut[49][9];
              muxOutConnector[25] = fifoOut[50][9];
              muxOutConnector[26] = fifoOut[17][2];
              muxOutConnector[27] = fifoOut[18][2];
              muxOutConnector[28] = fifoOut[19][2];
              muxOutConnector[29] = fifoOut[20][2];
              muxOutConnector[30] = fifoOut[21][2];
              muxOutConnector[31] = fifoOut[22][2];
              muxOutConnector[32] = fifoOut[23][2];
              muxOutConnector[33] = fifoOut[24][2];
              muxOutConnector[34] = fifoOut[25][2];
              muxOutConnector[35] = fifoOut[0][1];
              muxOutConnector[36] = fifoOut[1][1];
              muxOutConnector[37] = fifoOut[2][1];
              muxOutConnector[38] = fifoOut[3][1];
              muxOutConnector[39] = fifoOut[4][1];
              muxOutConnector[40] = fifoOut[5][1];
              muxOutConnector[41] = fifoOut[6][1];
              muxOutConnector[42] = fifoOut[7][1];
              muxOutConnector[43] = fifoOut[8][1];
              muxOutConnector[44] = fifoOut[9][1];
              muxOutConnector[45] = fifoOut[10][1];
              muxOutConnector[46] = fifoOut[11][1];
              muxOutConnector[47] = fifoOut[12][1];
              muxOutConnector[48] = fifoOut[13][1];
              muxOutConnector[49] = fifoOut[14][1];
              muxOutConnector[50] = fifoOut[15][1];
              muxOutConnector[51] = fifoOut[16][1];
       end
       17: begin
              muxOutConnector[0] = fifoOut[51][10];
              muxOutConnector[1] = fifoOut[26][9];
              muxOutConnector[2] = fifoOut[27][9];
              muxOutConnector[3] = fifoOut[28][9];
              muxOutConnector[4] = fifoOut[29][9];
              muxOutConnector[5] = fifoOut[30][9];
              muxOutConnector[6] = fifoOut[31][9];
              muxOutConnector[7] = fifoOut[32][9];
              muxOutConnector[8] = fifoOut[33][9];
              muxOutConnector[9] = fifoOut[34][9];
              muxOutConnector[10] = fifoOut[35][9];
              muxOutConnector[11] = fifoOut[36][9];
              muxOutConnector[12] = fifoOut[37][9];
              muxOutConnector[13] = fifoOut[38][9];
              muxOutConnector[14] = fifoOut[39][9];
              muxOutConnector[15] = fifoOut[40][9];
              muxOutConnector[16] = fifoOut[41][9];
              muxOutConnector[17] = fifoOut[42][9];
              muxOutConnector[18] = fifoOut[43][9];
              muxOutConnector[19] = fifoOut[44][9];
              muxOutConnector[20] = fifoOut[45][9];
              muxOutConnector[21] = fifoOut[46][9];
              muxOutConnector[22] = fifoOut[47][9];
              muxOutConnector[23] = fifoOut[48][9];
              muxOutConnector[24] = fifoOut[49][9];
              muxOutConnector[25] = fifoOut[50][9];
              muxOutConnector[26] = fifoOut[17][2];
              muxOutConnector[27] = fifoOut[18][2];
              muxOutConnector[28] = fifoOut[19][2];
              muxOutConnector[29] = fifoOut[20][2];
              muxOutConnector[30] = fifoOut[21][2];
              muxOutConnector[31] = fifoOut[22][2];
              muxOutConnector[32] = fifoOut[23][2];
              muxOutConnector[33] = fifoOut[24][2];
              muxOutConnector[34] = fifoOut[25][2];
              muxOutConnector[35] = fifoOut[0][1];
              muxOutConnector[36] = fifoOut[1][1];
              muxOutConnector[37] = fifoOut[2][1];
              muxOutConnector[38] = fifoOut[3][1];
              muxOutConnector[39] = fifoOut[4][1];
              muxOutConnector[40] = fifoOut[5][1];
              muxOutConnector[41] = fifoOut[6][1];
              muxOutConnector[42] = fifoOut[7][1];
              muxOutConnector[43] = fifoOut[8][1];
              muxOutConnector[44] = fifoOut[9][1];
              muxOutConnector[45] = fifoOut[10][1];
              muxOutConnector[46] = fifoOut[11][1];
              muxOutConnector[47] = fifoOut[12][1];
              muxOutConnector[48] = fifoOut[13][1];
              muxOutConnector[49] = fifoOut[14][1];
              muxOutConnector[50] = fifoOut[15][1];
              muxOutConnector[51] = fifoOut[16][1];
       end
       18: begin
              muxOutConnector[0] = fifoOut[51][10];
              muxOutConnector[1] = fifoOut[26][9];
              muxOutConnector[2] = fifoOut[27][9];
              muxOutConnector[3] = fifoOut[28][9];
              muxOutConnector[4] = fifoOut[29][9];
              muxOutConnector[5] = fifoOut[30][9];
              muxOutConnector[6] = fifoOut[31][9];
              muxOutConnector[7] = fifoOut[32][9];
              muxOutConnector[8] = fifoOut[33][9];
              muxOutConnector[9] = fifoOut[34][9];
              muxOutConnector[10] = fifoOut[35][9];
              muxOutConnector[11] = fifoOut[36][9];
              muxOutConnector[12] = fifoOut[37][9];
              muxOutConnector[13] = fifoOut[38][9];
              muxOutConnector[14] = fifoOut[39][9];
              muxOutConnector[15] = fifoOut[40][9];
              muxOutConnector[16] = fifoOut[41][9];
              muxOutConnector[17] = fifoOut[42][9];
              muxOutConnector[18] = fifoOut[43][9];
              muxOutConnector[19] = fifoOut[44][9];
              muxOutConnector[20] = fifoOut[45][9];
              muxOutConnector[21] = fifoOut[46][9];
              muxOutConnector[22] = fifoOut[47][9];
              muxOutConnector[23] = fifoOut[48][9];
              muxOutConnector[24] = fifoOut[49][9];
              muxOutConnector[25] = fifoOut[50][9];
              muxOutConnector[26] = fifoOut[17][2];
              muxOutConnector[27] = fifoOut[18][2];
              muxOutConnector[28] = fifoOut[19][2];
              muxOutConnector[29] = fifoOut[20][2];
              muxOutConnector[30] = fifoOut[21][2];
              muxOutConnector[31] = fifoOut[22][2];
              muxOutConnector[32] = fifoOut[23][2];
              muxOutConnector[33] = fifoOut[24][2];
              muxOutConnector[34] = fifoOut[25][2];
              muxOutConnector[35] = fifoOut[0][1];
              muxOutConnector[36] = fifoOut[1][1];
              muxOutConnector[37] = fifoOut[2][1];
              muxOutConnector[38] = fifoOut[3][1];
              muxOutConnector[39] = fifoOut[4][1];
              muxOutConnector[40] = fifoOut[5][1];
              muxOutConnector[41] = fifoOut[6][1];
              muxOutConnector[42] = fifoOut[7][1];
              muxOutConnector[43] = fifoOut[8][1];
              muxOutConnector[44] = fifoOut[9][1];
              muxOutConnector[45] = fifoOut[10][1];
              muxOutConnector[46] = fifoOut[11][1];
              muxOutConnector[47] = fifoOut[12][1];
              muxOutConnector[48] = fifoOut[13][1];
              muxOutConnector[49] = fifoOut[14][1];
              muxOutConnector[50] = fifoOut[15][1];
              muxOutConnector[51] = fifoOut[16][1];
       end
       19: begin
              muxOutConnector[0] = fifoOut[51][10];
              muxOutConnector[1] = fifoOut[26][9];
              muxOutConnector[2] = fifoOut[27][9];
              muxOutConnector[3] = fifoOut[28][9];
              muxOutConnector[4] = fifoOut[29][9];
              muxOutConnector[5] = fifoOut[30][9];
              muxOutConnector[6] = fifoOut[31][9];
              muxOutConnector[7] = fifoOut[32][9];
              muxOutConnector[8] = fifoOut[33][9];
              muxOutConnector[9] = fifoOut[34][9];
              muxOutConnector[10] = fifoOut[35][9];
              muxOutConnector[11] = fifoOut[36][9];
              muxOutConnector[12] = fifoOut[37][9];
              muxOutConnector[13] = fifoOut[38][9];
              muxOutConnector[14] = fifoOut[39][9];
              muxOutConnector[15] = fifoOut[40][9];
              muxOutConnector[16] = fifoOut[41][9];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[17][2];
              muxOutConnector[27] = fifoOut[18][2];
              muxOutConnector[28] = fifoOut[19][2];
              muxOutConnector[29] = fifoOut[20][2];
              muxOutConnector[30] = fifoOut[21][2];
              muxOutConnector[31] = fifoOut[22][2];
              muxOutConnector[32] = fifoOut[23][2];
              muxOutConnector[33] = fifoOut[24][2];
              muxOutConnector[34] = fifoOut[25][2];
              muxOutConnector[35] = fifoOut[0][1];
              muxOutConnector[36] = fifoOut[1][1];
              muxOutConnector[37] = fifoOut[2][1];
              muxOutConnector[38] = fifoOut[3][1];
              muxOutConnector[39] = fifoOut[4][1];
              muxOutConnector[40] = fifoOut[5][1];
              muxOutConnector[41] = fifoOut[6][1];
              muxOutConnector[42] = fifoOut[7][1];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
