`timescale 1ns / 1ps
module LMem0To1_511_circ12_ys_scripted(
        muxOut,
        ly0In,
        wr_en,
        feedback_en,
        rd_address,
        rd_en,
        clk,
        rst
);
input feedback_en;
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 16;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        if(feedback_en) begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= fifoOut[i][c-1];
         end
        end
        else begin
         for(i = r-1; i > -1; i=i-1) begin
              fifoOut[i][0] <= ly0InConnector[i];
         end
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[10][10];
              muxOutConnector[1] = fifoOut[11][10];
              muxOutConnector[2] = fifoOut[12][10];
              muxOutConnector[3] = fifoOut[13][10];
              muxOutConnector[4] = fifoOut[14][10];
              muxOutConnector[5] = fifoOut[15][10];
              muxOutConnector[6] = fifoOut[16][10];
              muxOutConnector[7] = fifoOut[17][10];
              muxOutConnector[8] = fifoOut[18][10];
              muxOutConnector[9] = fifoOut[19][10];
              muxOutConnector[10] = fifoOut[20][10];
              muxOutConnector[11] = fifoOut[21][10];
              muxOutConnector[12] = fifoOut[22][10];
              muxOutConnector[13] = fifoOut[23][10];
              muxOutConnector[14] = fifoOut[24][10];
              muxOutConnector[15] = fifoOut[25][10];
              muxOutConnector[16] = fifoOut[0][9];
              muxOutConnector[17] = fifoOut[1][9];
              muxOutConnector[18] = fifoOut[2][9];
              muxOutConnector[19] = fifoOut[3][9];
              muxOutConnector[20] = fifoOut[4][9];
              muxOutConnector[21] = fifoOut[5][9];
              muxOutConnector[22] = fifoOut[6][9];
              muxOutConnector[23] = fifoOut[7][9];
              muxOutConnector[24] = fifoOut[8][9];
              muxOutConnector[25] = fifoOut[9][9];
              muxOutConnector[26] = fifoOut[25][2];
              muxOutConnector[27] = fifoOut[0][1];
              muxOutConnector[28] = fifoOut[1][1];
              muxOutConnector[29] = fifoOut[2][1];
              muxOutConnector[30] = fifoOut[3][1];
              muxOutConnector[31] = fifoOut[4][1];
              muxOutConnector[32] = fifoOut[5][1];
              muxOutConnector[33] = fifoOut[6][1];
              muxOutConnector[34] = fifoOut[7][1];
              muxOutConnector[35] = fifoOut[8][1];
              muxOutConnector[36] = fifoOut[9][1];
              muxOutConnector[37] = fifoOut[10][1];
              muxOutConnector[38] = fifoOut[11][1];
              muxOutConnector[39] = fifoOut[12][1];
              muxOutConnector[40] = fifoOut[13][1];
              muxOutConnector[41] = fifoOut[14][1];
              muxOutConnector[42] = fifoOut[15][1];
              muxOutConnector[43] = fifoOut[16][1];
              muxOutConnector[44] = fifoOut[17][1];
              muxOutConnector[45] = fifoOut[18][1];
              muxOutConnector[46] = fifoOut[19][1];
              muxOutConnector[47] = fifoOut[20][1];
              muxOutConnector[48] = fifoOut[21][1];
              muxOutConnector[49] = fifoOut[22][1];
              muxOutConnector[50] = fifoOut[23][1];
              muxOutConnector[51] = fifoOut[24][1];
       end
       1: begin
              muxOutConnector[0] = fifoOut[10][10];
              muxOutConnector[1] = fifoOut[11][10];
              muxOutConnector[2] = fifoOut[12][10];
              muxOutConnector[3] = fifoOut[13][10];
              muxOutConnector[4] = fifoOut[14][10];
              muxOutConnector[5] = fifoOut[15][10];
              muxOutConnector[6] = fifoOut[16][10];
              muxOutConnector[7] = fifoOut[17][10];
              muxOutConnector[8] = fifoOut[18][10];
              muxOutConnector[9] = fifoOut[19][10];
              muxOutConnector[10] = fifoOut[20][10];
              muxOutConnector[11] = fifoOut[21][10];
              muxOutConnector[12] = fifoOut[22][10];
              muxOutConnector[13] = fifoOut[23][10];
              muxOutConnector[14] = fifoOut[24][10];
              muxOutConnector[15] = fifoOut[25][10];
              muxOutConnector[16] = fifoOut[0][9];
              muxOutConnector[17] = fifoOut[1][9];
              muxOutConnector[18] = fifoOut[2][9];
              muxOutConnector[19] = fifoOut[3][9];
              muxOutConnector[20] = fifoOut[4][9];
              muxOutConnector[21] = fifoOut[5][9];
              muxOutConnector[22] = fifoOut[6][9];
              muxOutConnector[23] = fifoOut[7][9];
              muxOutConnector[24] = fifoOut[8][9];
              muxOutConnector[25] = fifoOut[9][9];
              muxOutConnector[26] = fifoOut[25][2];
              muxOutConnector[27] = fifoOut[0][1];
              muxOutConnector[28] = fifoOut[1][1];
              muxOutConnector[29] = fifoOut[2][1];
              muxOutConnector[30] = fifoOut[3][1];
              muxOutConnector[31] = fifoOut[4][1];
              muxOutConnector[32] = fifoOut[5][1];
              muxOutConnector[33] = fifoOut[6][1];
              muxOutConnector[34] = fifoOut[7][1];
              muxOutConnector[35] = fifoOut[8][1];
              muxOutConnector[36] = fifoOut[9][1];
              muxOutConnector[37] = fifoOut[10][1];
              muxOutConnector[38] = fifoOut[11][1];
              muxOutConnector[39] = fifoOut[12][1];
              muxOutConnector[40] = fifoOut[13][1];
              muxOutConnector[41] = fifoOut[14][1];
              muxOutConnector[42] = fifoOut[15][1];
              muxOutConnector[43] = fifoOut[16][1];
              muxOutConnector[44] = fifoOut[34][0];
              muxOutConnector[45] = fifoOut[35][0];
              muxOutConnector[46] = fifoOut[36][0];
              muxOutConnector[47] = fifoOut[37][0];
              muxOutConnector[48] = fifoOut[38][0];
              muxOutConnector[49] = fifoOut[39][0];
              muxOutConnector[50] = fifoOut[40][0];
              muxOutConnector[51] = fifoOut[41][0];
       end
       2: begin
              muxOutConnector[0] = fifoOut[10][10];
              muxOutConnector[1] = fifoOut[11][10];
              muxOutConnector[2] = fifoOut[12][10];
              muxOutConnector[3] = fifoOut[13][10];
              muxOutConnector[4] = fifoOut[14][10];
              muxOutConnector[5] = fifoOut[15][10];
              muxOutConnector[6] = fifoOut[16][10];
              muxOutConnector[7] = fifoOut[17][10];
              muxOutConnector[8] = fifoOut[18][10];
              muxOutConnector[9] = fifoOut[19][10];
              muxOutConnector[10] = fifoOut[20][10];
              muxOutConnector[11] = fifoOut[21][10];
              muxOutConnector[12] = fifoOut[22][10];
              muxOutConnector[13] = fifoOut[23][10];
              muxOutConnector[14] = fifoOut[24][10];
              muxOutConnector[15] = fifoOut[25][10];
              muxOutConnector[16] = fifoOut[0][9];
              muxOutConnector[17] = fifoOut[1][9];
              muxOutConnector[18] = fifoOut[2][9];
              muxOutConnector[19] = fifoOut[3][9];
              muxOutConnector[20] = fifoOut[4][9];
              muxOutConnector[21] = fifoOut[5][9];
              muxOutConnector[22] = fifoOut[6][9];
              muxOutConnector[23] = fifoOut[7][9];
              muxOutConnector[24] = fifoOut[8][9];
              muxOutConnector[25] = fifoOut[9][9];
              muxOutConnector[26] = fifoOut[42][1];
              muxOutConnector[27] = fifoOut[43][1];
              muxOutConnector[28] = fifoOut[44][1];
              muxOutConnector[29] = fifoOut[45][1];
              muxOutConnector[30] = fifoOut[46][1];
              muxOutConnector[31] = fifoOut[47][1];
              muxOutConnector[32] = fifoOut[48][1];
              muxOutConnector[33] = fifoOut[49][1];
              muxOutConnector[34] = fifoOut[50][1];
              muxOutConnector[35] = fifoOut[51][1];
              muxOutConnector[36] = fifoOut[26][0];
              muxOutConnector[37] = fifoOut[27][0];
              muxOutConnector[38] = fifoOut[28][0];
              muxOutConnector[39] = fifoOut[29][0];
              muxOutConnector[40] = fifoOut[30][0];
              muxOutConnector[41] = fifoOut[31][0];
              muxOutConnector[42] = fifoOut[32][0];
              muxOutConnector[43] = fifoOut[33][0];
              muxOutConnector[44] = fifoOut[34][0];
              muxOutConnector[45] = fifoOut[35][0];
              muxOutConnector[46] = fifoOut[36][0];
              muxOutConnector[47] = fifoOut[37][0];
              muxOutConnector[48] = fifoOut[38][0];
              muxOutConnector[49] = fifoOut[39][0];
              muxOutConnector[50] = fifoOut[40][0];
              muxOutConnector[51] = fifoOut[41][0];
       end
       3: begin
              muxOutConnector[0] = fifoOut[10][10];
              muxOutConnector[1] = fifoOut[11][10];
              muxOutConnector[2] = fifoOut[12][10];
              muxOutConnector[3] = fifoOut[13][10];
              muxOutConnector[4] = fifoOut[14][10];
              muxOutConnector[5] = fifoOut[15][10];
              muxOutConnector[6] = fifoOut[16][10];
              muxOutConnector[7] = fifoOut[17][10];
              muxOutConnector[8] = fifoOut[18][10];
              muxOutConnector[9] = fifoOut[19][10];
              muxOutConnector[10] = fifoOut[20][10];
              muxOutConnector[11] = fifoOut[21][10];
              muxOutConnector[12] = fifoOut[22][10];
              muxOutConnector[13] = fifoOut[23][10];
              muxOutConnector[14] = fifoOut[24][10];
              muxOutConnector[15] = fifoOut[25][10];
              muxOutConnector[16] = fifoOut[0][9];
              muxOutConnector[17] = fifoOut[1][9];
              muxOutConnector[18] = fifoOut[2][9];
              muxOutConnector[19] = fifoOut[3][9];
              muxOutConnector[20] = fifoOut[4][9];
              muxOutConnector[21] = fifoOut[5][9];
              muxOutConnector[22] = fifoOut[6][9];
              muxOutConnector[23] = fifoOut[7][9];
              muxOutConnector[24] = fifoOut[8][9];
              muxOutConnector[25] = fifoOut[9][9];
              muxOutConnector[26] = fifoOut[42][1];
              muxOutConnector[27] = fifoOut[43][1];
              muxOutConnector[28] = fifoOut[44][1];
              muxOutConnector[29] = fifoOut[45][1];
              muxOutConnector[30] = fifoOut[46][1];
              muxOutConnector[31] = fifoOut[47][1];
              muxOutConnector[32] = fifoOut[48][1];
              muxOutConnector[33] = fifoOut[49][1];
              muxOutConnector[34] = fifoOut[50][1];
              muxOutConnector[35] = fifoOut[51][1];
              muxOutConnector[36] = fifoOut[26][0];
              muxOutConnector[37] = fifoOut[27][0];
              muxOutConnector[38] = fifoOut[28][0];
              muxOutConnector[39] = fifoOut[29][0];
              muxOutConnector[40] = fifoOut[30][0];
              muxOutConnector[41] = fifoOut[31][0];
              muxOutConnector[42] = fifoOut[32][0];
              muxOutConnector[43] = fifoOut[33][0];
              muxOutConnector[44] = fifoOut[34][0];
              muxOutConnector[45] = fifoOut[35][0];
              muxOutConnector[46] = fifoOut[36][0];
              muxOutConnector[47] = fifoOut[37][0];
              muxOutConnector[48] = fifoOut[38][0];
              muxOutConnector[49] = fifoOut[39][0];
              muxOutConnector[50] = fifoOut[40][0];
              muxOutConnector[51] = fifoOut[41][0];
       end
       4: begin
              muxOutConnector[0] = fifoOut[10][10];
              muxOutConnector[1] = fifoOut[11][10];
              muxOutConnector[2] = fifoOut[12][10];
              muxOutConnector[3] = fifoOut[13][10];
              muxOutConnector[4] = fifoOut[14][10];
              muxOutConnector[5] = fifoOut[15][10];
              muxOutConnector[6] = fifoOut[16][10];
              muxOutConnector[7] = fifoOut[17][10];
              muxOutConnector[8] = fifoOut[18][10];
              muxOutConnector[9] = fifoOut[19][10];
              muxOutConnector[10] = fifoOut[20][10];
              muxOutConnector[11] = fifoOut[21][10];
              muxOutConnector[12] = fifoOut[22][10];
              muxOutConnector[13] = fifoOut[23][10];
              muxOutConnector[14] = fifoOut[24][10];
              muxOutConnector[15] = fifoOut[25][10];
              muxOutConnector[16] = fifoOut[0][9];
              muxOutConnector[17] = fifoOut[1][9];
              muxOutConnector[18] = fifoOut[2][9];
              muxOutConnector[19] = fifoOut[3][9];
              muxOutConnector[20] = fifoOut[4][9];
              muxOutConnector[21] = fifoOut[5][9];
              muxOutConnector[22] = fifoOut[6][9];
              muxOutConnector[23] = fifoOut[7][9];
              muxOutConnector[24] = fifoOut[8][9];
              muxOutConnector[25] = fifoOut[9][9];
              muxOutConnector[26] = fifoOut[42][1];
              muxOutConnector[27] = fifoOut[43][1];
              muxOutConnector[28] = fifoOut[44][1];
              muxOutConnector[29] = fifoOut[45][1];
              muxOutConnector[30] = fifoOut[46][1];
              muxOutConnector[31] = fifoOut[47][1];
              muxOutConnector[32] = fifoOut[48][1];
              muxOutConnector[33] = fifoOut[49][1];
              muxOutConnector[34] = fifoOut[50][1];
              muxOutConnector[35] = fifoOut[51][1];
              muxOutConnector[36] = fifoOut[26][0];
              muxOutConnector[37] = fifoOut[27][0];
              muxOutConnector[38] = fifoOut[28][0];
              muxOutConnector[39] = fifoOut[29][0];
              muxOutConnector[40] = fifoOut[30][0];
              muxOutConnector[41] = fifoOut[31][0];
              muxOutConnector[42] = fifoOut[32][0];
              muxOutConnector[43] = fifoOut[33][0];
              muxOutConnector[44] = fifoOut[34][0];
              muxOutConnector[45] = fifoOut[35][0];
              muxOutConnector[46] = fifoOut[36][0];
              muxOutConnector[47] = fifoOut[37][0];
              muxOutConnector[48] = fifoOut[38][0];
              muxOutConnector[49] = fifoOut[39][0];
              muxOutConnector[50] = fifoOut[40][0];
              muxOutConnector[51] = fifoOut[41][0];
       end
       5: begin
              muxOutConnector[0] = fifoOut[10][10];
              muxOutConnector[1] = fifoOut[11][10];
              muxOutConnector[2] = fifoOut[12][10];
              muxOutConnector[3] = fifoOut[13][10];
              muxOutConnector[4] = fifoOut[14][10];
              muxOutConnector[5] = fifoOut[15][10];
              muxOutConnector[6] = fifoOut[16][10];
              muxOutConnector[7] = fifoOut[17][10];
              muxOutConnector[8] = fifoOut[18][10];
              muxOutConnector[9] = fifoOut[19][10];
              muxOutConnector[10] = fifoOut[20][10];
              muxOutConnector[11] = fifoOut[21][10];
              muxOutConnector[12] = fifoOut[22][10];
              muxOutConnector[13] = fifoOut[23][10];
              muxOutConnector[14] = fifoOut[24][10];
              muxOutConnector[15] = fifoOut[25][10];
              muxOutConnector[16] = fifoOut[0][9];
              muxOutConnector[17] = fifoOut[1][9];
              muxOutConnector[18] = fifoOut[2][9];
              muxOutConnector[19] = fifoOut[3][9];
              muxOutConnector[20] = fifoOut[4][9];
              muxOutConnector[21] = fifoOut[5][9];
              muxOutConnector[22] = fifoOut[6][9];
              muxOutConnector[23] = fifoOut[7][9];
              muxOutConnector[24] = fifoOut[8][9];
              muxOutConnector[25] = fifoOut[9][9];
              muxOutConnector[26] = fifoOut[42][1];
              muxOutConnector[27] = fifoOut[43][1];
              muxOutConnector[28] = fifoOut[44][1];
              muxOutConnector[29] = fifoOut[45][1];
              muxOutConnector[30] = fifoOut[46][1];
              muxOutConnector[31] = fifoOut[47][1];
              muxOutConnector[32] = fifoOut[48][1];
              muxOutConnector[33] = fifoOut[49][1];
              muxOutConnector[34] = fifoOut[50][1];
              muxOutConnector[35] = fifoOut[51][1];
              muxOutConnector[36] = fifoOut[26][0];
              muxOutConnector[37] = fifoOut[27][0];
              muxOutConnector[38] = fifoOut[28][0];
              muxOutConnector[39] = fifoOut[29][0];
              muxOutConnector[40] = fifoOut[30][0];
              muxOutConnector[41] = fifoOut[31][0];
              muxOutConnector[42] = fifoOut[32][0];
              muxOutConnector[43] = fifoOut[33][0];
              muxOutConnector[44] = fifoOut[0][4];
              muxOutConnector[45] = fifoOut[1][4];
              muxOutConnector[46] = fifoOut[2][4];
              muxOutConnector[47] = fifoOut[3][4];
              muxOutConnector[48] = fifoOut[4][4];
              muxOutConnector[49] = fifoOut[5][4];
              muxOutConnector[50] = fifoOut[6][4];
              muxOutConnector[51] = fifoOut[7][4];
       end
       6: begin
              muxOutConnector[0] = fifoOut[10][10];
              muxOutConnector[1] = fifoOut[11][10];
              muxOutConnector[2] = fifoOut[12][10];
              muxOutConnector[3] = fifoOut[13][10];
              muxOutConnector[4] = fifoOut[14][10];
              muxOutConnector[5] = fifoOut[15][10];
              muxOutConnector[6] = fifoOut[16][10];
              muxOutConnector[7] = fifoOut[17][10];
              muxOutConnector[8] = fifoOut[18][10];
              muxOutConnector[9] = fifoOut[19][10];
              muxOutConnector[10] = fifoOut[20][10];
              muxOutConnector[11] = fifoOut[21][10];
              muxOutConnector[12] = fifoOut[22][10];
              muxOutConnector[13] = fifoOut[23][10];
              muxOutConnector[14] = fifoOut[24][10];
              muxOutConnector[15] = fifoOut[25][10];
              muxOutConnector[16] = fifoOut[0][9];
              muxOutConnector[17] = fifoOut[1][9];
              muxOutConnector[18] = fifoOut[2][9];
              muxOutConnector[19] = fifoOut[3][9];
              muxOutConnector[20] = fifoOut[4][9];
              muxOutConnector[21] = fifoOut[5][9];
              muxOutConnector[22] = fifoOut[6][9];
              muxOutConnector[23] = fifoOut[7][9];
              muxOutConnector[24] = fifoOut[8][9];
              muxOutConnector[25] = fifoOut[9][9];
              muxOutConnector[26] = fifoOut[8][5];
              muxOutConnector[27] = fifoOut[9][5];
              muxOutConnector[28] = fifoOut[10][5];
              muxOutConnector[29] = fifoOut[11][5];
              muxOutConnector[30] = fifoOut[12][5];
              muxOutConnector[31] = fifoOut[13][5];
              muxOutConnector[32] = fifoOut[14][5];
              muxOutConnector[33] = fifoOut[15][5];
              muxOutConnector[34] = fifoOut[16][5];
              muxOutConnector[35] = fifoOut[17][5];
              muxOutConnector[36] = fifoOut[18][5];
              muxOutConnector[37] = fifoOut[19][5];
              muxOutConnector[38] = fifoOut[20][5];
              muxOutConnector[39] = fifoOut[21][5];
              muxOutConnector[40] = fifoOut[22][5];
              muxOutConnector[41] = fifoOut[23][5];
              muxOutConnector[42] = fifoOut[24][5];
              muxOutConnector[43] = fifoOut[25][5];
              muxOutConnector[44] = fifoOut[0][4];
              muxOutConnector[45] = fifoOut[1][4];
              muxOutConnector[46] = fifoOut[2][4];
              muxOutConnector[47] = fifoOut[3][4];
              muxOutConnector[48] = fifoOut[4][4];
              muxOutConnector[49] = fifoOut[5][4];
              muxOutConnector[50] = fifoOut[6][4];
              muxOutConnector[51] = fifoOut[7][4];
       end
       7: begin
              muxOutConnector[0] = fifoOut[10][10];
              muxOutConnector[1] = fifoOut[11][10];
              muxOutConnector[2] = fifoOut[12][10];
              muxOutConnector[3] = fifoOut[13][10];
              muxOutConnector[4] = fifoOut[14][10];
              muxOutConnector[5] = fifoOut[15][10];
              muxOutConnector[6] = fifoOut[16][10];
              muxOutConnector[7] = fifoOut[17][10];
              muxOutConnector[8] = fifoOut[18][10];
              muxOutConnector[9] = fifoOut[19][10];
              muxOutConnector[10] = fifoOut[20][10];
              muxOutConnector[11] = fifoOut[21][10];
              muxOutConnector[12] = fifoOut[22][10];
              muxOutConnector[13] = fifoOut[23][10];
              muxOutConnector[14] = fifoOut[24][10];
              muxOutConnector[15] = fifoOut[25][10];
              muxOutConnector[16] = fifoOut[0][9];
              muxOutConnector[17] = fifoOut[1][9];
              muxOutConnector[18] = fifoOut[2][9];
              muxOutConnector[19] = fifoOut[3][9];
              muxOutConnector[20] = fifoOut[4][9];
              muxOutConnector[21] = fifoOut[5][9];
              muxOutConnector[22] = fifoOut[6][9];
              muxOutConnector[23] = fifoOut[7][9];
              muxOutConnector[24] = fifoOut[8][9];
              muxOutConnector[25] = fifoOut[9][9];
              muxOutConnector[26] = fifoOut[8][5];
              muxOutConnector[27] = fifoOut[9][5];
              muxOutConnector[28] = fifoOut[10][5];
              muxOutConnector[29] = fifoOut[11][5];
              muxOutConnector[30] = fifoOut[12][5];
              muxOutConnector[31] = fifoOut[13][5];
              muxOutConnector[32] = fifoOut[14][5];
              muxOutConnector[33] = fifoOut[15][5];
              muxOutConnector[34] = fifoOut[16][5];
              muxOutConnector[35] = fifoOut[17][5];
              muxOutConnector[36] = fifoOut[18][5];
              muxOutConnector[37] = fifoOut[19][5];
              muxOutConnector[38] = fifoOut[20][5];
              muxOutConnector[39] = fifoOut[21][5];
              muxOutConnector[40] = fifoOut[22][5];
              muxOutConnector[41] = fifoOut[23][5];
              muxOutConnector[42] = fifoOut[24][5];
              muxOutConnector[43] = fifoOut[25][5];
              muxOutConnector[44] = fifoOut[0][4];
              muxOutConnector[45] = fifoOut[1][4];
              muxOutConnector[46] = fifoOut[2][4];
              muxOutConnector[47] = fifoOut[3][4];
              muxOutConnector[48] = fifoOut[4][4];
              muxOutConnector[49] = fifoOut[5][4];
              muxOutConnector[50] = fifoOut[6][4];
              muxOutConnector[51] = fifoOut[7][4];
       end
       8: begin
              muxOutConnector[0] = fifoOut[10][10];
              muxOutConnector[1] = fifoOut[11][10];
              muxOutConnector[2] = fifoOut[12][10];
              muxOutConnector[3] = fifoOut[13][10];
              muxOutConnector[4] = fifoOut[14][10];
              muxOutConnector[5] = fifoOut[15][10];
              muxOutConnector[6] = fifoOut[16][10];
              muxOutConnector[7] = fifoOut[17][10];
              muxOutConnector[8] = fifoOut[18][10];
              muxOutConnector[9] = fifoOut[19][10];
              muxOutConnector[10] = fifoOut[20][10];
              muxOutConnector[11] = fifoOut[21][10];
              muxOutConnector[12] = fifoOut[22][10];
              muxOutConnector[13] = fifoOut[23][10];
              muxOutConnector[14] = fifoOut[24][10];
              muxOutConnector[15] = fifoOut[25][10];
              muxOutConnector[16] = fifoOut[0][9];
              muxOutConnector[17] = fifoOut[1][9];
              muxOutConnector[18] = fifoOut[2][9];
              muxOutConnector[19] = fifoOut[3][9];
              muxOutConnector[20] = fifoOut[4][9];
              muxOutConnector[21] = fifoOut[5][9];
              muxOutConnector[22] = fifoOut[6][9];
              muxOutConnector[23] = fifoOut[7][9];
              muxOutConnector[24] = fifoOut[8][9];
              muxOutConnector[25] = fifoOut[9][9];
              muxOutConnector[26] = fifoOut[8][5];
              muxOutConnector[27] = fifoOut[9][5];
              muxOutConnector[28] = fifoOut[10][5];
              muxOutConnector[29] = fifoOut[11][5];
              muxOutConnector[30] = fifoOut[12][5];
              muxOutConnector[31] = fifoOut[13][5];
              muxOutConnector[32] = fifoOut[14][5];
              muxOutConnector[33] = fifoOut[15][5];
              muxOutConnector[34] = fifoOut[16][5];
              muxOutConnector[35] = fifoOut[17][5];
              muxOutConnector[36] = fifoOut[18][5];
              muxOutConnector[37] = fifoOut[19][5];
              muxOutConnector[38] = fifoOut[20][5];
              muxOutConnector[39] = fifoOut[21][5];
              muxOutConnector[40] = fifoOut[22][5];
              muxOutConnector[41] = fifoOut[23][5];
              muxOutConnector[42] = fifoOut[24][5];
              muxOutConnector[43] = fifoOut[25][5];
              muxOutConnector[44] = fifoOut[0][4];
              muxOutConnector[45] = fifoOut[1][4];
              muxOutConnector[46] = fifoOut[2][4];
              muxOutConnector[47] = fifoOut[3][4];
              muxOutConnector[48] = fifoOut[4][4];
              muxOutConnector[49] = fifoOut[5][4];
              muxOutConnector[50] = fifoOut[6][4];
              muxOutConnector[51] = fifoOut[7][4];
       end
       9: begin
              muxOutConnector[0] = fifoOut[10][10];
              muxOutConnector[1] = fifoOut[11][10];
              muxOutConnector[2] = fifoOut[12][10];
              muxOutConnector[3] = fifoOut[13][10];
              muxOutConnector[4] = fifoOut[14][10];
              muxOutConnector[5] = fifoOut[15][10];
              muxOutConnector[6] = fifoOut[16][10];
              muxOutConnector[7] = fifoOut[17][10];
              muxOutConnector[8] = fifoOut[18][10];
              muxOutConnector[9] = fifoOut[19][10];
              muxOutConnector[10] = fifoOut[20][10];
              muxOutConnector[11] = fifoOut[21][10];
              muxOutConnector[12] = fifoOut[22][10];
              muxOutConnector[13] = fifoOut[23][10];
              muxOutConnector[14] = fifoOut[24][10];
              muxOutConnector[15] = fifoOut[25][10];
              muxOutConnector[16] = fifoOut[0][9];
              muxOutConnector[17] = fifoOut[1][9];
              muxOutConnector[18] = fifoOut[2][9];
              muxOutConnector[19] = fifoOut[3][9];
              muxOutConnector[20] = fifoOut[4][9];
              muxOutConnector[21] = fifoOut[5][9];
              muxOutConnector[22] = fifoOut[6][9];
              muxOutConnector[23] = fifoOut[7][9];
              muxOutConnector[24] = fifoOut[8][9];
              muxOutConnector[25] = fifoOut[9][9];
              muxOutConnector[26] = fifoOut[8][5];
              muxOutConnector[27] = fifoOut[9][5];
              muxOutConnector[28] = fifoOut[10][5];
              muxOutConnector[29] = fifoOut[11][5];
              muxOutConnector[30] = fifoOut[12][5];
              muxOutConnector[31] = fifoOut[13][5];
              muxOutConnector[32] = fifoOut[14][5];
              muxOutConnector[33] = fifoOut[15][5];
              muxOutConnector[34] = fifoOut[16][5];
              muxOutConnector[35] = fifoOut[17][5];
              muxOutConnector[36] = fifoOut[18][5];
              muxOutConnector[37] = fifoOut[19][5];
              muxOutConnector[38] = fifoOut[20][5];
              muxOutConnector[39] = fifoOut[21][5];
              muxOutConnector[40] = fifoOut[22][5];
              muxOutConnector[41] = fifoOut[23][5];
              muxOutConnector[42] = fifoOut[24][5];
              muxOutConnector[43] = fifoOut[25][5];
              muxOutConnector[44] = fifoOut[0][4];
              muxOutConnector[45] = fifoOut[1][4];
              muxOutConnector[46] = fifoOut[2][4];
              muxOutConnector[47] = fifoOut[3][4];
              muxOutConnector[48] = fifoOut[4][4];
              muxOutConnector[49] = fifoOut[5][4];
              muxOutConnector[50] = fifoOut[6][4];
              muxOutConnector[51] = fifoOut[7][4];
       end
       10: begin
              muxOutConnector[0] = fifoOut[10][10];
              muxOutConnector[1] = fifoOut[11][10];
              muxOutConnector[2] = fifoOut[12][10];
              muxOutConnector[3] = fifoOut[13][10];
              muxOutConnector[4] = fifoOut[14][10];
              muxOutConnector[5] = fifoOut[15][10];
              muxOutConnector[6] = fifoOut[16][10];
              muxOutConnector[7] = fifoOut[34][9];
              muxOutConnector[8] = fifoOut[35][9];
              muxOutConnector[9] = fifoOut[36][9];
              muxOutConnector[10] = fifoOut[37][9];
              muxOutConnector[11] = fifoOut[38][9];
              muxOutConnector[12] = fifoOut[39][9];
              muxOutConnector[13] = fifoOut[40][9];
              muxOutConnector[14] = fifoOut[41][9];
              muxOutConnector[15] = fifoOut[42][9];
              muxOutConnector[16] = fifoOut[43][9];
              muxOutConnector[17] = fifoOut[44][9];
              muxOutConnector[18] = fifoOut[45][9];
              muxOutConnector[19] = fifoOut[46][9];
              muxOutConnector[20] = fifoOut[47][9];
              muxOutConnector[21] = fifoOut[48][9];
              muxOutConnector[22] = fifoOut[49][9];
              muxOutConnector[23] = fifoOut[50][9];
              muxOutConnector[24] = fifoOut[51][9];
              muxOutConnector[25] = fifoOut[26][8];
              muxOutConnector[26] = fifoOut[8][5];
              muxOutConnector[27] = fifoOut[9][5];
              muxOutConnector[28] = fifoOut[10][5];
              muxOutConnector[29] = fifoOut[11][5];
              muxOutConnector[30] = fifoOut[12][5];
              muxOutConnector[31] = fifoOut[13][5];
              muxOutConnector[32] = fifoOut[14][5];
              muxOutConnector[33] = fifoOut[15][5];
              muxOutConnector[34] = fifoOut[16][5];
              muxOutConnector[35] = fifoOut[17][5];
              muxOutConnector[36] = fifoOut[18][5];
              muxOutConnector[37] = fifoOut[19][5];
              muxOutConnector[38] = fifoOut[20][5];
              muxOutConnector[39] = fifoOut[21][5];
              muxOutConnector[40] = fifoOut[22][5];
              muxOutConnector[41] = fifoOut[23][5];
              muxOutConnector[42] = fifoOut[24][5];
              muxOutConnector[43] = fifoOut[25][5];
              muxOutConnector[44] = fifoOut[0][4];
              muxOutConnector[45] = fifoOut[1][4];
              muxOutConnector[46] = fifoOut[2][4];
              muxOutConnector[47] = fifoOut[3][4];
              muxOutConnector[48] = fifoOut[4][4];
              muxOutConnector[49] = fifoOut[5][4];
              muxOutConnector[50] = fifoOut[6][4];
              muxOutConnector[51] = fifoOut[7][4];
       end
       11: begin
              muxOutConnector[0] = fifoOut[27][9];
              muxOutConnector[1] = fifoOut[28][9];
              muxOutConnector[2] = fifoOut[29][9];
              muxOutConnector[3] = fifoOut[30][9];
              muxOutConnector[4] = fifoOut[31][9];
              muxOutConnector[5] = fifoOut[32][9];
              muxOutConnector[6] = fifoOut[33][9];
              muxOutConnector[7] = fifoOut[34][9];
              muxOutConnector[8] = fifoOut[35][9];
              muxOutConnector[9] = fifoOut[36][9];
              muxOutConnector[10] = fifoOut[37][9];
              muxOutConnector[11] = fifoOut[38][9];
              muxOutConnector[12] = fifoOut[39][9];
              muxOutConnector[13] = fifoOut[40][9];
              muxOutConnector[14] = fifoOut[41][9];
              muxOutConnector[15] = fifoOut[42][9];
              muxOutConnector[16] = fifoOut[43][9];
              muxOutConnector[17] = fifoOut[44][9];
              muxOutConnector[18] = fifoOut[45][9];
              muxOutConnector[19] = fifoOut[46][9];
              muxOutConnector[20] = fifoOut[47][9];
              muxOutConnector[21] = fifoOut[48][9];
              muxOutConnector[22] = fifoOut[49][9];
              muxOutConnector[23] = fifoOut[50][9];
              muxOutConnector[24] = fifoOut[51][9];
              muxOutConnector[25] = fifoOut[26][8];
              muxOutConnector[26] = fifoOut[8][5];
              muxOutConnector[27] = fifoOut[9][5];
              muxOutConnector[28] = fifoOut[10][5];
              muxOutConnector[29] = fifoOut[11][5];
              muxOutConnector[30] = fifoOut[12][5];
              muxOutConnector[31] = fifoOut[13][5];
              muxOutConnector[32] = fifoOut[14][5];
              muxOutConnector[33] = fifoOut[15][5];
              muxOutConnector[34] = fifoOut[16][5];
              muxOutConnector[35] = fifoOut[17][5];
              muxOutConnector[36] = fifoOut[18][5];
              muxOutConnector[37] = fifoOut[19][5];
              muxOutConnector[38] = fifoOut[20][5];
              muxOutConnector[39] = fifoOut[21][5];
              muxOutConnector[40] = fifoOut[22][5];
              muxOutConnector[41] = fifoOut[23][5];
              muxOutConnector[42] = fifoOut[24][5];
              muxOutConnector[43] = fifoOut[25][5];
              muxOutConnector[44] = fifoOut[0][4];
              muxOutConnector[45] = fifoOut[1][4];
              muxOutConnector[46] = fifoOut[2][4];
              muxOutConnector[47] = fifoOut[3][4];
              muxOutConnector[48] = fifoOut[4][4];
              muxOutConnector[49] = fifoOut[5][4];
              muxOutConnector[50] = fifoOut[6][4];
              muxOutConnector[51] = fifoOut[7][4];
       end
       12: begin
              muxOutConnector[0] = fifoOut[27][9];
              muxOutConnector[1] = fifoOut[28][9];
              muxOutConnector[2] = fifoOut[29][9];
              muxOutConnector[3] = fifoOut[30][9];
              muxOutConnector[4] = fifoOut[31][9];
              muxOutConnector[5] = fifoOut[32][9];
              muxOutConnector[6] = fifoOut[33][9];
              muxOutConnector[7] = fifoOut[34][9];
              muxOutConnector[8] = fifoOut[35][9];
              muxOutConnector[9] = fifoOut[36][9];
              muxOutConnector[10] = fifoOut[37][9];
              muxOutConnector[11] = fifoOut[38][9];
              muxOutConnector[12] = fifoOut[39][9];
              muxOutConnector[13] = fifoOut[40][9];
              muxOutConnector[14] = fifoOut[41][9];
              muxOutConnector[15] = fifoOut[42][9];
              muxOutConnector[16] = fifoOut[43][9];
              muxOutConnector[17] = fifoOut[44][9];
              muxOutConnector[18] = fifoOut[45][9];
              muxOutConnector[19] = fifoOut[46][9];
              muxOutConnector[20] = fifoOut[47][9];
              muxOutConnector[21] = fifoOut[48][9];
              muxOutConnector[22] = fifoOut[49][9];
              muxOutConnector[23] = fifoOut[50][9];
              muxOutConnector[24] = fifoOut[51][9];
              muxOutConnector[25] = fifoOut[26][8];
              muxOutConnector[26] = fifoOut[8][5];
              muxOutConnector[27] = fifoOut[9][5];
              muxOutConnector[28] = fifoOut[10][5];
              muxOutConnector[29] = fifoOut[11][5];
              muxOutConnector[30] = fifoOut[12][5];
              muxOutConnector[31] = fifoOut[13][5];
              muxOutConnector[32] = fifoOut[14][5];
              muxOutConnector[33] = fifoOut[15][5];
              muxOutConnector[34] = fifoOut[16][5];
              muxOutConnector[35] = fifoOut[17][5];
              muxOutConnector[36] = fifoOut[18][5];
              muxOutConnector[37] = fifoOut[19][5];
              muxOutConnector[38] = fifoOut[20][5];
              muxOutConnector[39] = fifoOut[21][5];
              muxOutConnector[40] = fifoOut[22][5];
              muxOutConnector[41] = fifoOut[23][5];
              muxOutConnector[42] = fifoOut[24][5];
              muxOutConnector[43] = fifoOut[25][5];
              muxOutConnector[44] = fifoOut[0][4];
              muxOutConnector[45] = fifoOut[1][4];
              muxOutConnector[46] = fifoOut[2][4];
              muxOutConnector[47] = fifoOut[3][4];
              muxOutConnector[48] = fifoOut[4][4];
              muxOutConnector[49] = fifoOut[5][4];
              muxOutConnector[50] = fifoOut[6][4];
              muxOutConnector[51] = fifoOut[7][4];
       end
       13: begin
              muxOutConnector[0] = fifoOut[27][9];
              muxOutConnector[1] = fifoOut[28][9];
              muxOutConnector[2] = fifoOut[29][9];
              muxOutConnector[3] = fifoOut[30][9];
              muxOutConnector[4] = fifoOut[31][9];
              muxOutConnector[5] = fifoOut[32][9];
              muxOutConnector[6] = fifoOut[33][9];
              muxOutConnector[7] = fifoOut[34][9];
              muxOutConnector[8] = fifoOut[35][9];
              muxOutConnector[9] = fifoOut[36][9];
              muxOutConnector[10] = fifoOut[37][9];
              muxOutConnector[11] = fifoOut[38][9];
              muxOutConnector[12] = fifoOut[39][9];
              muxOutConnector[13] = fifoOut[40][9];
              muxOutConnector[14] = fifoOut[41][9];
              muxOutConnector[15] = fifoOut[42][9];
              muxOutConnector[16] = fifoOut[43][9];
              muxOutConnector[17] = fifoOut[44][9];
              muxOutConnector[18] = fifoOut[45][9];
              muxOutConnector[19] = fifoOut[46][9];
              muxOutConnector[20] = fifoOut[47][9];
              muxOutConnector[21] = fifoOut[48][9];
              muxOutConnector[22] = fifoOut[49][9];
              muxOutConnector[23] = fifoOut[50][9];
              muxOutConnector[24] = fifoOut[51][9];
              muxOutConnector[25] = fifoOut[26][8];
              muxOutConnector[26] = fifoOut[8][5];
              muxOutConnector[27] = fifoOut[9][5];
              muxOutConnector[28] = fifoOut[10][5];
              muxOutConnector[29] = fifoOut[11][5];
              muxOutConnector[30] = fifoOut[12][5];
              muxOutConnector[31] = fifoOut[13][5];
              muxOutConnector[32] = fifoOut[14][5];
              muxOutConnector[33] = fifoOut[15][5];
              muxOutConnector[34] = fifoOut[16][5];
              muxOutConnector[35] = fifoOut[17][5];
              muxOutConnector[36] = fifoOut[18][5];
              muxOutConnector[37] = fifoOut[19][5];
              muxOutConnector[38] = fifoOut[20][5];
              muxOutConnector[39] = fifoOut[21][5];
              muxOutConnector[40] = fifoOut[22][5];
              muxOutConnector[41] = fifoOut[23][5];
              muxOutConnector[42] = fifoOut[24][5];
              muxOutConnector[43] = fifoOut[25][5];
              muxOutConnector[44] = fifoOut[0][4];
              muxOutConnector[45] = fifoOut[1][4];
              muxOutConnector[46] = fifoOut[2][4];
              muxOutConnector[47] = fifoOut[3][4];
              muxOutConnector[48] = fifoOut[4][4];
              muxOutConnector[49] = fifoOut[5][4];
              muxOutConnector[50] = fifoOut[6][4];
              muxOutConnector[51] = fifoOut[7][4];
       end
       14: begin
              muxOutConnector[0] = fifoOut[27][9];
              muxOutConnector[1] = fifoOut[28][9];
              muxOutConnector[2] = fifoOut[29][9];
              muxOutConnector[3] = fifoOut[30][9];
              muxOutConnector[4] = fifoOut[31][9];
              muxOutConnector[5] = fifoOut[32][9];
              muxOutConnector[6] = fifoOut[33][9];
              muxOutConnector[7] = fifoOut[0][13];
              muxOutConnector[8] = fifoOut[1][13];
              muxOutConnector[9] = fifoOut[2][13];
              muxOutConnector[10] = fifoOut[3][13];
              muxOutConnector[11] = fifoOut[4][13];
              muxOutConnector[12] = fifoOut[5][13];
              muxOutConnector[13] = fifoOut[6][13];
              muxOutConnector[14] = fifoOut[7][13];
              muxOutConnector[15] = fifoOut[8][13];
              muxOutConnector[16] = fifoOut[9][13];
              muxOutConnector[17] = fifoOut[10][13];
              muxOutConnector[18] = fifoOut[11][13];
              muxOutConnector[19] = fifoOut[12][13];
              muxOutConnector[20] = fifoOut[13][13];
              muxOutConnector[21] = fifoOut[14][13];
              muxOutConnector[22] = fifoOut[15][13];
              muxOutConnector[23] = fifoOut[16][13];
              muxOutConnector[24] = fifoOut[17][13];
              muxOutConnector[25] = fifoOut[18][13];
              muxOutConnector[26] = fifoOut[8][5];
              muxOutConnector[27] = fifoOut[9][5];
              muxOutConnector[28] = fifoOut[10][5];
              muxOutConnector[29] = fifoOut[11][5];
              muxOutConnector[30] = fifoOut[12][5];
              muxOutConnector[31] = fifoOut[13][5];
              muxOutConnector[32] = fifoOut[14][5];
              muxOutConnector[33] = fifoOut[15][5];
              muxOutConnector[34] = fifoOut[16][5];
              muxOutConnector[35] = fifoOut[17][5];
              muxOutConnector[36] = fifoOut[18][5];
              muxOutConnector[37] = fifoOut[19][5];
              muxOutConnector[38] = fifoOut[20][5];
              muxOutConnector[39] = fifoOut[21][5];
              muxOutConnector[40] = fifoOut[22][5];
              muxOutConnector[41] = fifoOut[23][5];
              muxOutConnector[42] = fifoOut[24][5];
              muxOutConnector[43] = fifoOut[25][5];
              muxOutConnector[44] = fifoOut[0][4];
              muxOutConnector[45] = fifoOut[1][4];
              muxOutConnector[46] = fifoOut[2][4];
              muxOutConnector[47] = fifoOut[3][4];
              muxOutConnector[48] = fifoOut[4][4];
              muxOutConnector[49] = fifoOut[5][4];
              muxOutConnector[50] = fifoOut[6][4];
              muxOutConnector[51] = fifoOut[7][4];
       end
       15: begin
              muxOutConnector[0] = fifoOut[19][14];
              muxOutConnector[1] = fifoOut[20][14];
              muxOutConnector[2] = fifoOut[21][14];
              muxOutConnector[3] = fifoOut[22][14];
              muxOutConnector[4] = fifoOut[23][14];
              muxOutConnector[5] = fifoOut[24][14];
              muxOutConnector[6] = fifoOut[25][14];
              muxOutConnector[7] = fifoOut[0][13];
              muxOutConnector[8] = fifoOut[1][13];
              muxOutConnector[9] = fifoOut[2][13];
              muxOutConnector[10] = fifoOut[3][13];
              muxOutConnector[11] = fifoOut[4][13];
              muxOutConnector[12] = fifoOut[5][13];
              muxOutConnector[13] = fifoOut[6][13];
              muxOutConnector[14] = fifoOut[7][13];
              muxOutConnector[15] = fifoOut[8][13];
              muxOutConnector[16] = fifoOut[9][13];
              muxOutConnector[17] = fifoOut[10][13];
              muxOutConnector[18] = fifoOut[11][13];
              muxOutConnector[19] = fifoOut[12][13];
              muxOutConnector[20] = fifoOut[13][13];
              muxOutConnector[21] = fifoOut[14][13];
              muxOutConnector[22] = fifoOut[15][13];
              muxOutConnector[23] = fifoOut[16][13];
              muxOutConnector[24] = fifoOut[17][13];
              muxOutConnector[25] = fifoOut[18][13];
              muxOutConnector[26] = fifoOut[8][5];
              muxOutConnector[27] = fifoOut[9][5];
              muxOutConnector[28] = fifoOut[10][5];
              muxOutConnector[29] = fifoOut[11][5];
              muxOutConnector[30] = fifoOut[12][5];
              muxOutConnector[31] = fifoOut[13][5];
              muxOutConnector[32] = fifoOut[14][5];
              muxOutConnector[33] = fifoOut[15][5];
              muxOutConnector[34] = fifoOut[16][5];
              muxOutConnector[35] = fifoOut[17][5];
              muxOutConnector[36] = fifoOut[18][5];
              muxOutConnector[37] = fifoOut[19][5];
              muxOutConnector[38] = fifoOut[20][5];
              muxOutConnector[39] = fifoOut[21][5];
              muxOutConnector[40] = fifoOut[22][5];
              muxOutConnector[41] = fifoOut[23][5];
              muxOutConnector[42] = fifoOut[24][5];
              muxOutConnector[43] = fifoOut[25][5];
              muxOutConnector[44] = fifoOut[0][4];
              muxOutConnector[45] = fifoOut[1][4];
              muxOutConnector[46] = fifoOut[2][4];
              muxOutConnector[47] = fifoOut[3][4];
              muxOutConnector[48] = fifoOut[4][4];
              muxOutConnector[49] = fifoOut[5][4];
              muxOutConnector[50] = fifoOut[6][4];
              muxOutConnector[51] = fifoOut[7][4];
       end
       16: begin
              muxOutConnector[0] = fifoOut[19][14];
              muxOutConnector[1] = fifoOut[20][14];
              muxOutConnector[2] = fifoOut[21][14];
              muxOutConnector[3] = fifoOut[22][14];
              muxOutConnector[4] = fifoOut[23][14];
              muxOutConnector[5] = fifoOut[24][14];
              muxOutConnector[6] = fifoOut[25][14];
              muxOutConnector[7] = fifoOut[0][13];
              muxOutConnector[8] = fifoOut[1][13];
              muxOutConnector[9] = fifoOut[2][13];
              muxOutConnector[10] = fifoOut[3][13];
              muxOutConnector[11] = fifoOut[4][13];
              muxOutConnector[12] = fifoOut[5][13];
              muxOutConnector[13] = fifoOut[6][13];
              muxOutConnector[14] = fifoOut[7][13];
              muxOutConnector[15] = fifoOut[8][13];
              muxOutConnector[16] = fifoOut[9][13];
              muxOutConnector[17] = fifoOut[10][13];
              muxOutConnector[18] = fifoOut[11][13];
              muxOutConnector[19] = fifoOut[12][13];
              muxOutConnector[20] = fifoOut[13][13];
              muxOutConnector[21] = fifoOut[14][13];
              muxOutConnector[22] = fifoOut[15][13];
              muxOutConnector[23] = fifoOut[16][13];
              muxOutConnector[24] = fifoOut[17][13];
              muxOutConnector[25] = fifoOut[18][13];
              muxOutConnector[26] = fifoOut[8][5];
              muxOutConnector[27] = fifoOut[9][5];
              muxOutConnector[28] = fifoOut[10][5];
              muxOutConnector[29] = fifoOut[11][5];
              muxOutConnector[30] = fifoOut[12][5];
              muxOutConnector[31] = fifoOut[13][5];
              muxOutConnector[32] = fifoOut[14][5];
              muxOutConnector[33] = fifoOut[15][5];
              muxOutConnector[34] = fifoOut[16][5];
              muxOutConnector[35] = fifoOut[17][5];
              muxOutConnector[36] = fifoOut[18][5];
              muxOutConnector[37] = fifoOut[19][5];
              muxOutConnector[38] = fifoOut[20][5];
              muxOutConnector[39] = fifoOut[21][5];
              muxOutConnector[40] = fifoOut[22][5];
              muxOutConnector[41] = fifoOut[23][5];
              muxOutConnector[42] = fifoOut[24][5];
              muxOutConnector[43] = fifoOut[25][5];
              muxOutConnector[44] = fifoOut[0][4];
              muxOutConnector[45] = fifoOut[1][4];
              muxOutConnector[46] = fifoOut[2][4];
              muxOutConnector[47] = fifoOut[3][4];
              muxOutConnector[48] = fifoOut[4][4];
              muxOutConnector[49] = fifoOut[5][4];
              muxOutConnector[50] = fifoOut[6][4];
              muxOutConnector[51] = fifoOut[7][4];
       end
       17: begin
              muxOutConnector[0] = fifoOut[19][14];
              muxOutConnector[1] = fifoOut[20][14];
              muxOutConnector[2] = fifoOut[21][14];
              muxOutConnector[3] = fifoOut[22][14];
              muxOutConnector[4] = fifoOut[23][14];
              muxOutConnector[5] = fifoOut[24][14];
              muxOutConnector[6] = fifoOut[25][14];
              muxOutConnector[7] = fifoOut[0][13];
              muxOutConnector[8] = fifoOut[1][13];
              muxOutConnector[9] = fifoOut[2][13];
              muxOutConnector[10] = fifoOut[3][13];
              muxOutConnector[11] = fifoOut[4][13];
              muxOutConnector[12] = fifoOut[5][13];
              muxOutConnector[13] = fifoOut[6][13];
              muxOutConnector[14] = fifoOut[7][13];
              muxOutConnector[15] = fifoOut[8][13];
              muxOutConnector[16] = fifoOut[9][13];
              muxOutConnector[17] = fifoOut[10][13];
              muxOutConnector[18] = fifoOut[11][13];
              muxOutConnector[19] = fifoOut[12][13];
              muxOutConnector[20] = fifoOut[13][13];
              muxOutConnector[21] = fifoOut[14][13];
              muxOutConnector[22] = fifoOut[15][13];
              muxOutConnector[23] = fifoOut[16][13];
              muxOutConnector[24] = fifoOut[17][13];
              muxOutConnector[25] = fifoOut[18][13];
              muxOutConnector[26] = fifoOut[8][5];
              muxOutConnector[27] = fifoOut[9][5];
              muxOutConnector[28] = fifoOut[10][5];
              muxOutConnector[29] = fifoOut[11][5];
              muxOutConnector[30] = fifoOut[12][5];
              muxOutConnector[31] = fifoOut[13][5];
              muxOutConnector[32] = fifoOut[14][5];
              muxOutConnector[33] = fifoOut[15][5];
              muxOutConnector[34] = fifoOut[16][5];
              muxOutConnector[35] = fifoOut[17][5];
              muxOutConnector[36] = fifoOut[18][5];
              muxOutConnector[37] = fifoOut[19][5];
              muxOutConnector[38] = fifoOut[20][5];
              muxOutConnector[39] = fifoOut[21][5];
              muxOutConnector[40] = fifoOut[22][5];
              muxOutConnector[41] = fifoOut[23][5];
              muxOutConnector[42] = fifoOut[24][5];
              muxOutConnector[43] = fifoOut[25][5];
              muxOutConnector[44] = fifoOut[0][4];
              muxOutConnector[45] = fifoOut[1][4];
              muxOutConnector[46] = fifoOut[2][4];
              muxOutConnector[47] = fifoOut[3][4];
              muxOutConnector[48] = fifoOut[4][4];
              muxOutConnector[49] = fifoOut[5][4];
              muxOutConnector[50] = fifoOut[6][4];
              muxOutConnector[51] = fifoOut[7][4];
       end
       18: begin
              muxOutConnector[0] = fifoOut[19][14];
              muxOutConnector[1] = fifoOut[20][14];
              muxOutConnector[2] = fifoOut[21][14];
              muxOutConnector[3] = fifoOut[22][14];
              muxOutConnector[4] = fifoOut[23][14];
              muxOutConnector[5] = fifoOut[24][14];
              muxOutConnector[6] = fifoOut[25][14];
              muxOutConnector[7] = fifoOut[0][13];
              muxOutConnector[8] = fifoOut[1][13];
              muxOutConnector[9] = fifoOut[2][13];
              muxOutConnector[10] = fifoOut[3][13];
              muxOutConnector[11] = fifoOut[4][13];
              muxOutConnector[12] = fifoOut[5][13];
              muxOutConnector[13] = fifoOut[6][13];
              muxOutConnector[14] = fifoOut[7][13];
              muxOutConnector[15] = fifoOut[8][13];
              muxOutConnector[16] = fifoOut[9][13];
              muxOutConnector[17] = fifoOut[10][13];
              muxOutConnector[18] = fifoOut[11][13];
              muxOutConnector[19] = fifoOut[12][13];
              muxOutConnector[20] = fifoOut[13][13];
              muxOutConnector[21] = fifoOut[14][13];
              muxOutConnector[22] = fifoOut[15][13];
              muxOutConnector[23] = fifoOut[16][13];
              muxOutConnector[24] = fifoOut[17][13];
              muxOutConnector[25] = fifoOut[18][13];
              muxOutConnector[26] = fifoOut[8][5];
              muxOutConnector[27] = fifoOut[9][5];
              muxOutConnector[28] = fifoOut[10][5];
              muxOutConnector[29] = fifoOut[11][5];
              muxOutConnector[30] = fifoOut[12][5];
              muxOutConnector[31] = fifoOut[13][5];
              muxOutConnector[32] = fifoOut[14][5];
              muxOutConnector[33] = fifoOut[15][5];
              muxOutConnector[34] = fifoOut[16][5];
              muxOutConnector[35] = fifoOut[17][5];
              muxOutConnector[36] = fifoOut[18][5];
              muxOutConnector[37] = fifoOut[19][5];
              muxOutConnector[38] = fifoOut[20][5];
              muxOutConnector[39] = fifoOut[21][5];
              muxOutConnector[40] = fifoOut[22][5];
              muxOutConnector[41] = fifoOut[23][5];
              muxOutConnector[42] = fifoOut[24][5];
              muxOutConnector[43] = fifoOut[25][5];
              muxOutConnector[44] = fifoOut[0][4];
              muxOutConnector[45] = fifoOut[1][4];
              muxOutConnector[46] = fifoOut[2][4];
              muxOutConnector[47] = fifoOut[3][4];
              muxOutConnector[48] = fifoOut[4][4];
              muxOutConnector[49] = fifoOut[5][4];
              muxOutConnector[50] = fifoOut[6][4];
              muxOutConnector[51] = fifoOut[7][4];
       end
       19: begin
              muxOutConnector[0] = fifoOut[19][14];
              muxOutConnector[1] = fifoOut[20][14];
              muxOutConnector[2] = fifoOut[21][14];
              muxOutConnector[3] = fifoOut[22][14];
              muxOutConnector[4] = fifoOut[23][14];
              muxOutConnector[5] = fifoOut[24][14];
              muxOutConnector[6] = fifoOut[25][14];
              muxOutConnector[7] = fifoOut[0][13];
              muxOutConnector[8] = fifoOut[1][13];
              muxOutConnector[9] = fifoOut[2][13];
              muxOutConnector[10] = fifoOut[3][13];
              muxOutConnector[11] = fifoOut[4][13];
              muxOutConnector[12] = fifoOut[5][13];
              muxOutConnector[13] = fifoOut[6][13];
              muxOutConnector[14] = fifoOut[7][13];
              muxOutConnector[15] = fifoOut[8][13];
              muxOutConnector[16] = fifoOut[9][13];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[8][5];
              muxOutConnector[27] = fifoOut[9][5];
              muxOutConnector[28] = fifoOut[10][5];
              muxOutConnector[29] = fifoOut[11][5];
              muxOutConnector[30] = fifoOut[12][5];
              muxOutConnector[31] = fifoOut[13][5];
              muxOutConnector[32] = fifoOut[14][5];
              muxOutConnector[33] = fifoOut[15][5];
              muxOutConnector[34] = fifoOut[16][5];
              muxOutConnector[35] = fifoOut[17][5];
              muxOutConnector[36] = fifoOut[18][5];
              muxOutConnector[37] = fifoOut[19][5];
              muxOutConnector[38] = fifoOut[20][5];
              muxOutConnector[39] = fifoOut[21][5];
              muxOutConnector[40] = fifoOut[22][5];
              muxOutConnector[41] = fifoOut[23][5];
              muxOutConnector[42] = fifoOut[24][5];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
