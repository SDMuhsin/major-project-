`timescale 1ns / 1ps
module LMem0To1_511_circ8_ys_scripted(
        muxOut,
        ly0In,
        wr_en,
        rd_address,
        rd_en,
        clk,
        rst
);
parameter w = 6; // DataWidth
parameter r = 52;
parameter c = 13;
parameter ADDRESSWIDTH = 5;
parameter muxOutSymbols = 52;
parameter maxVal = 6'b011111;
parameter READDISABLEDCASE = 5'd31; // if rd_en is 0 go to a default Address 

output [ muxOutSymbols * w - 1 : 0]muxOut;
input [ r * w - 1 : 0 ]ly0In; // Change #3
input wr_en;
input [ADDRESSWIDTH-1:0]rd_address;
input rd_en;
input clk,rst; // #C

wire [ADDRESSWIDTH-1:0]rd_address_case;
wire [w-1:0]ly0InConnector[r-1:0]; // Change #
reg [w-1:0]muxOutConnector[ muxOutSymbols  - 1 : 0];
reg [w-1:0] fifoOut[r-1:0][c-1:0]; // FIFO Outputs

genvar k;
generate
    for (k=0;k<muxOutSymbols;k=k+1)begin:assign_output
        assign muxOut[ (k+1)*w-1:k*w] = muxOutConnector[k];
    end
endgenerate
generate
    for (k=0;k<r;k=k+1)begin:assign_input
        assign ly0InConnector[k] = ly0In[(k+1)*w-1:k*w];
    end
endgenerate

integer i;
integer j;

always@(posedge clk)begin
    if (rst) begin
        for(i=0;i<r;i=i+1)begin
            for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= 0;
            end
        end
    end
    else if(wr_en) begin
        // Shift
        for(i = r-1; i > -1; i=i-1) begin
            for(j= c-1; j > 0; j=j-1)begin
                fifoOut[i][j] <=  fifoOut[i][j-1];
            end
        end
        // Input
        for(i = r-1; i > -1; i=i-1) begin
            fifoOut[i][0] <= ly0InConnector[i];
        end
    end
    else begin
        for(i=0;i<r;i=i+1)begin
           for(j=0;j<c;j=j+1)begin
                fifoOut[i][j] <= fifoOut[i][j];
           end
        end
    end
end

assign rd_address_case = rd_en ? rd_address : READDISABLEDCASE;

always@(*)begin
    case(rd_address_case)
       0: begin
              muxOutConnector[0] = fifoOut[13][9];
              muxOutConnector[1] = fifoOut[14][9];
              muxOutConnector[2] = fifoOut[15][9];
              muxOutConnector[3] = fifoOut[16][9];
              muxOutConnector[4] = fifoOut[17][9];
              muxOutConnector[5] = fifoOut[18][9];
              muxOutConnector[6] = fifoOut[19][9];
              muxOutConnector[7] = fifoOut[20][9];
              muxOutConnector[8] = fifoOut[21][9];
              muxOutConnector[9] = fifoOut[22][9];
              muxOutConnector[10] = fifoOut[23][9];
              muxOutConnector[11] = fifoOut[24][9];
              muxOutConnector[12] = fifoOut[25][9];
              muxOutConnector[13] = fifoOut[0][8];
              muxOutConnector[14] = fifoOut[1][8];
              muxOutConnector[15] = fifoOut[2][8];
              muxOutConnector[16] = fifoOut[3][8];
              muxOutConnector[17] = fifoOut[4][8];
              muxOutConnector[18] = fifoOut[5][8];
              muxOutConnector[19] = fifoOut[6][8];
              muxOutConnector[20] = fifoOut[7][8];
              muxOutConnector[21] = fifoOut[8][8];
              muxOutConnector[22] = fifoOut[9][8];
              muxOutConnector[23] = fifoOut[10][8];
              muxOutConnector[24] = fifoOut[11][8];
              muxOutConnector[25] = fifoOut[12][8];
              muxOutConnector[26] = fifoOut[14][3];
              muxOutConnector[27] = fifoOut[15][3];
              muxOutConnector[28] = fifoOut[16][3];
              muxOutConnector[29] = fifoOut[17][3];
              muxOutConnector[30] = fifoOut[18][3];
              muxOutConnector[31] = fifoOut[19][3];
              muxOutConnector[32] = fifoOut[20][3];
              muxOutConnector[33] = fifoOut[21][3];
              muxOutConnector[34] = fifoOut[22][3];
              muxOutConnector[35] = fifoOut[23][3];
              muxOutConnector[36] = fifoOut[24][3];
              muxOutConnector[37] = fifoOut[25][3];
              muxOutConnector[38] = fifoOut[0][2];
              muxOutConnector[39] = fifoOut[1][2];
              muxOutConnector[40] = fifoOut[2][2];
              muxOutConnector[41] = fifoOut[3][2];
              muxOutConnector[42] = fifoOut[4][2];
              muxOutConnector[43] = fifoOut[5][2];
              muxOutConnector[44] = fifoOut[6][2];
              muxOutConnector[45] = fifoOut[7][2];
              muxOutConnector[46] = fifoOut[8][2];
              muxOutConnector[47] = fifoOut[9][2];
              muxOutConnector[48] = fifoOut[10][2];
              muxOutConnector[49] = fifoOut[11][2];
              muxOutConnector[50] = fifoOut[12][2];
              muxOutConnector[51] = fifoOut[13][2];
       end
       1: begin
              muxOutConnector[0] = fifoOut[13][9];
              muxOutConnector[1] = fifoOut[14][9];
              muxOutConnector[2] = fifoOut[15][9];
              muxOutConnector[3] = fifoOut[16][9];
              muxOutConnector[4] = fifoOut[17][9];
              muxOutConnector[5] = fifoOut[18][9];
              muxOutConnector[6] = fifoOut[19][9];
              muxOutConnector[7] = fifoOut[20][9];
              muxOutConnector[8] = fifoOut[21][9];
              muxOutConnector[9] = fifoOut[22][9];
              muxOutConnector[10] = fifoOut[23][9];
              muxOutConnector[11] = fifoOut[24][9];
              muxOutConnector[12] = fifoOut[25][9];
              muxOutConnector[13] = fifoOut[0][8];
              muxOutConnector[14] = fifoOut[1][8];
              muxOutConnector[15] = fifoOut[2][8];
              muxOutConnector[16] = fifoOut[3][8];
              muxOutConnector[17] = fifoOut[4][8];
              muxOutConnector[18] = fifoOut[5][8];
              muxOutConnector[19] = fifoOut[6][8];
              muxOutConnector[20] = fifoOut[7][8];
              muxOutConnector[21] = fifoOut[8][8];
              muxOutConnector[22] = fifoOut[9][8];
              muxOutConnector[23] = fifoOut[10][8];
              muxOutConnector[24] = fifoOut[11][8];
              muxOutConnector[25] = fifoOut[12][8];
              muxOutConnector[26] = fifoOut[14][3];
              muxOutConnector[27] = fifoOut[15][3];
              muxOutConnector[28] = fifoOut[16][3];
              muxOutConnector[29] = fifoOut[17][3];
              muxOutConnector[30] = fifoOut[18][3];
              muxOutConnector[31] = fifoOut[19][3];
              muxOutConnector[32] = fifoOut[20][3];
              muxOutConnector[33] = fifoOut[21][3];
              muxOutConnector[34] = fifoOut[22][3];
              muxOutConnector[35] = fifoOut[23][3];
              muxOutConnector[36] = fifoOut[24][3];
              muxOutConnector[37] = fifoOut[25][3];
              muxOutConnector[38] = fifoOut[0][2];
              muxOutConnector[39] = fifoOut[1][2];
              muxOutConnector[40] = fifoOut[2][2];
              muxOutConnector[41] = fifoOut[3][2];
              muxOutConnector[42] = fifoOut[4][2];
              muxOutConnector[43] = fifoOut[5][2];
              muxOutConnector[44] = fifoOut[6][2];
              muxOutConnector[45] = fifoOut[7][2];
              muxOutConnector[46] = fifoOut[8][2];
              muxOutConnector[47] = fifoOut[9][2];
              muxOutConnector[48] = fifoOut[10][2];
              muxOutConnector[49] = fifoOut[11][2];
              muxOutConnector[50] = fifoOut[12][2];
              muxOutConnector[51] = fifoOut[13][2];
       end
       2: begin
              muxOutConnector[0] = fifoOut[13][9];
              muxOutConnector[1] = fifoOut[14][9];
              muxOutConnector[2] = fifoOut[15][9];
              muxOutConnector[3] = fifoOut[16][9];
              muxOutConnector[4] = fifoOut[17][9];
              muxOutConnector[5] = fifoOut[18][9];
              muxOutConnector[6] = fifoOut[19][9];
              muxOutConnector[7] = fifoOut[20][9];
              muxOutConnector[8] = fifoOut[21][9];
              muxOutConnector[9] = fifoOut[22][9];
              muxOutConnector[10] = fifoOut[23][9];
              muxOutConnector[11] = fifoOut[24][9];
              muxOutConnector[12] = fifoOut[25][9];
              muxOutConnector[13] = fifoOut[0][8];
              muxOutConnector[14] = fifoOut[1][8];
              muxOutConnector[15] = fifoOut[2][8];
              muxOutConnector[16] = fifoOut[3][8];
              muxOutConnector[17] = fifoOut[4][8];
              muxOutConnector[18] = fifoOut[5][8];
              muxOutConnector[19] = fifoOut[6][8];
              muxOutConnector[20] = fifoOut[7][8];
              muxOutConnector[21] = fifoOut[8][8];
              muxOutConnector[22] = fifoOut[9][8];
              muxOutConnector[23] = fifoOut[10][8];
              muxOutConnector[24] = fifoOut[11][8];
              muxOutConnector[25] = fifoOut[12][8];
              muxOutConnector[26] = fifoOut[14][3];
              muxOutConnector[27] = fifoOut[15][3];
              muxOutConnector[28] = fifoOut[16][3];
              muxOutConnector[29] = fifoOut[17][3];
              muxOutConnector[30] = fifoOut[18][3];
              muxOutConnector[31] = fifoOut[19][3];
              muxOutConnector[32] = fifoOut[20][3];
              muxOutConnector[33] = fifoOut[21][3];
              muxOutConnector[34] = fifoOut[22][3];
              muxOutConnector[35] = fifoOut[23][3];
              muxOutConnector[36] = fifoOut[24][3];
              muxOutConnector[37] = fifoOut[25][3];
              muxOutConnector[38] = fifoOut[0][2];
              muxOutConnector[39] = fifoOut[1][2];
              muxOutConnector[40] = fifoOut[2][2];
              muxOutConnector[41] = fifoOut[3][2];
              muxOutConnector[42] = fifoOut[4][2];
              muxOutConnector[43] = fifoOut[5][2];
              muxOutConnector[44] = fifoOut[6][2];
              muxOutConnector[45] = fifoOut[7][2];
              muxOutConnector[46] = fifoOut[8][2];
              muxOutConnector[47] = fifoOut[9][2];
              muxOutConnector[48] = fifoOut[10][2];
              muxOutConnector[49] = fifoOut[11][2];
              muxOutConnector[50] = fifoOut[12][2];
              muxOutConnector[51] = fifoOut[13][2];
       end
       3: begin
              muxOutConnector[0] = fifoOut[13][9];
              muxOutConnector[1] = fifoOut[14][9];
              muxOutConnector[2] = fifoOut[15][9];
              muxOutConnector[3] = fifoOut[16][9];
              muxOutConnector[4] = fifoOut[17][9];
              muxOutConnector[5] = fifoOut[18][9];
              muxOutConnector[6] = fifoOut[19][9];
              muxOutConnector[7] = fifoOut[20][9];
              muxOutConnector[8] = fifoOut[21][9];
              muxOutConnector[9] = fifoOut[22][9];
              muxOutConnector[10] = fifoOut[23][9];
              muxOutConnector[11] = fifoOut[24][9];
              muxOutConnector[12] = fifoOut[25][9];
              muxOutConnector[13] = fifoOut[0][8];
              muxOutConnector[14] = fifoOut[1][8];
              muxOutConnector[15] = fifoOut[2][8];
              muxOutConnector[16] = fifoOut[3][8];
              muxOutConnector[17] = fifoOut[4][8];
              muxOutConnector[18] = fifoOut[5][8];
              muxOutConnector[19] = fifoOut[6][8];
              muxOutConnector[20] = fifoOut[7][8];
              muxOutConnector[21] = fifoOut[8][8];
              muxOutConnector[22] = fifoOut[9][8];
              muxOutConnector[23] = fifoOut[10][8];
              muxOutConnector[24] = fifoOut[11][8];
              muxOutConnector[25] = fifoOut[12][8];
              muxOutConnector[26] = fifoOut[14][3];
              muxOutConnector[27] = fifoOut[15][3];
              muxOutConnector[28] = fifoOut[16][3];
              muxOutConnector[29] = fifoOut[48][2];
              muxOutConnector[30] = fifoOut[49][2];
              muxOutConnector[31] = fifoOut[50][2];
              muxOutConnector[32] = fifoOut[51][2];
              muxOutConnector[33] = fifoOut[26][1];
              muxOutConnector[34] = fifoOut[27][1];
              muxOutConnector[35] = fifoOut[28][1];
              muxOutConnector[36] = fifoOut[29][1];
              muxOutConnector[37] = fifoOut[30][1];
              muxOutConnector[38] = fifoOut[31][1];
              muxOutConnector[39] = fifoOut[32][1];
              muxOutConnector[40] = fifoOut[33][1];
              muxOutConnector[41] = fifoOut[34][1];
              muxOutConnector[42] = fifoOut[35][1];
              muxOutConnector[43] = fifoOut[36][1];
              muxOutConnector[44] = fifoOut[37][1];
              muxOutConnector[45] = fifoOut[38][1];
              muxOutConnector[46] = fifoOut[39][1];
              muxOutConnector[47] = fifoOut[40][1];
              muxOutConnector[48] = fifoOut[41][1];
              muxOutConnector[49] = fifoOut[42][1];
              muxOutConnector[50] = fifoOut[43][1];
              muxOutConnector[51] = fifoOut[44][1];
       end
       4: begin
              muxOutConnector[0] = fifoOut[13][9];
              muxOutConnector[1] = fifoOut[14][9];
              muxOutConnector[2] = fifoOut[15][9];
              muxOutConnector[3] = fifoOut[16][9];
              muxOutConnector[4] = fifoOut[17][9];
              muxOutConnector[5] = fifoOut[18][9];
              muxOutConnector[6] = fifoOut[19][9];
              muxOutConnector[7] = fifoOut[20][9];
              muxOutConnector[8] = fifoOut[21][9];
              muxOutConnector[9] = fifoOut[22][9];
              muxOutConnector[10] = fifoOut[23][9];
              muxOutConnector[11] = fifoOut[24][9];
              muxOutConnector[12] = fifoOut[25][9];
              muxOutConnector[13] = fifoOut[0][8];
              muxOutConnector[14] = fifoOut[1][8];
              muxOutConnector[15] = fifoOut[2][8];
              muxOutConnector[16] = fifoOut[3][8];
              muxOutConnector[17] = fifoOut[4][8];
              muxOutConnector[18] = fifoOut[5][8];
              muxOutConnector[19] = fifoOut[6][8];
              muxOutConnector[20] = fifoOut[7][8];
              muxOutConnector[21] = fifoOut[8][8];
              muxOutConnector[22] = fifoOut[9][8];
              muxOutConnector[23] = fifoOut[10][8];
              muxOutConnector[24] = fifoOut[11][8];
              muxOutConnector[25] = fifoOut[12][8];
              muxOutConnector[26] = fifoOut[45][2];
              muxOutConnector[27] = fifoOut[46][2];
              muxOutConnector[28] = fifoOut[47][2];
              muxOutConnector[29] = fifoOut[48][2];
              muxOutConnector[30] = fifoOut[49][2];
              muxOutConnector[31] = fifoOut[50][2];
              muxOutConnector[32] = fifoOut[51][2];
              muxOutConnector[33] = fifoOut[26][1];
              muxOutConnector[34] = fifoOut[27][1];
              muxOutConnector[35] = fifoOut[28][1];
              muxOutConnector[36] = fifoOut[29][1];
              muxOutConnector[37] = fifoOut[30][1];
              muxOutConnector[38] = fifoOut[31][1];
              muxOutConnector[39] = fifoOut[32][1];
              muxOutConnector[40] = fifoOut[33][1];
              muxOutConnector[41] = fifoOut[34][1];
              muxOutConnector[42] = fifoOut[35][1];
              muxOutConnector[43] = fifoOut[36][1];
              muxOutConnector[44] = fifoOut[37][1];
              muxOutConnector[45] = fifoOut[38][1];
              muxOutConnector[46] = fifoOut[39][1];
              muxOutConnector[47] = fifoOut[40][1];
              muxOutConnector[48] = fifoOut[41][1];
              muxOutConnector[49] = fifoOut[42][1];
              muxOutConnector[50] = fifoOut[43][1];
              muxOutConnector[51] = fifoOut[44][1];
       end
       5: begin
              muxOutConnector[0] = fifoOut[13][9];
              muxOutConnector[1] = fifoOut[14][9];
              muxOutConnector[2] = fifoOut[15][9];
              muxOutConnector[3] = fifoOut[16][9];
              muxOutConnector[4] = fifoOut[17][9];
              muxOutConnector[5] = fifoOut[18][9];
              muxOutConnector[6] = fifoOut[19][9];
              muxOutConnector[7] = fifoOut[20][9];
              muxOutConnector[8] = fifoOut[21][9];
              muxOutConnector[9] = fifoOut[22][9];
              muxOutConnector[10] = fifoOut[23][9];
              muxOutConnector[11] = fifoOut[24][9];
              muxOutConnector[12] = fifoOut[25][9];
              muxOutConnector[13] = fifoOut[0][8];
              muxOutConnector[14] = fifoOut[1][8];
              muxOutConnector[15] = fifoOut[2][8];
              muxOutConnector[16] = fifoOut[3][8];
              muxOutConnector[17] = fifoOut[4][8];
              muxOutConnector[18] = fifoOut[5][8];
              muxOutConnector[19] = fifoOut[6][8];
              muxOutConnector[20] = fifoOut[7][8];
              muxOutConnector[21] = fifoOut[8][8];
              muxOutConnector[22] = fifoOut[9][8];
              muxOutConnector[23] = fifoOut[10][8];
              muxOutConnector[24] = fifoOut[11][8];
              muxOutConnector[25] = fifoOut[12][8];
              muxOutConnector[26] = fifoOut[45][2];
              muxOutConnector[27] = fifoOut[46][2];
              muxOutConnector[28] = fifoOut[47][2];
              muxOutConnector[29] = fifoOut[48][2];
              muxOutConnector[30] = fifoOut[49][2];
              muxOutConnector[31] = fifoOut[50][2];
              muxOutConnector[32] = fifoOut[51][2];
              muxOutConnector[33] = fifoOut[26][1];
              muxOutConnector[34] = fifoOut[27][1];
              muxOutConnector[35] = fifoOut[28][1];
              muxOutConnector[36] = fifoOut[29][1];
              muxOutConnector[37] = fifoOut[30][1];
              muxOutConnector[38] = fifoOut[31][1];
              muxOutConnector[39] = fifoOut[32][1];
              muxOutConnector[40] = fifoOut[33][1];
              muxOutConnector[41] = fifoOut[34][1];
              muxOutConnector[42] = fifoOut[35][1];
              muxOutConnector[43] = fifoOut[36][1];
              muxOutConnector[44] = fifoOut[37][1];
              muxOutConnector[45] = fifoOut[38][1];
              muxOutConnector[46] = fifoOut[39][1];
              muxOutConnector[47] = fifoOut[40][1];
              muxOutConnector[48] = fifoOut[41][1];
              muxOutConnector[49] = fifoOut[42][1];
              muxOutConnector[50] = fifoOut[43][1];
              muxOutConnector[51] = fifoOut[44][1];
       end
       6: begin
              muxOutConnector[0] = fifoOut[13][9];
              muxOutConnector[1] = fifoOut[14][9];
              muxOutConnector[2] = fifoOut[15][9];
              muxOutConnector[3] = fifoOut[16][9];
              muxOutConnector[4] = fifoOut[17][9];
              muxOutConnector[5] = fifoOut[18][9];
              muxOutConnector[6] = fifoOut[19][9];
              muxOutConnector[7] = fifoOut[20][9];
              muxOutConnector[8] = fifoOut[21][9];
              muxOutConnector[9] = fifoOut[22][9];
              muxOutConnector[10] = fifoOut[23][9];
              muxOutConnector[11] = fifoOut[24][9];
              muxOutConnector[12] = fifoOut[25][9];
              muxOutConnector[13] = fifoOut[0][8];
              muxOutConnector[14] = fifoOut[1][8];
              muxOutConnector[15] = fifoOut[2][8];
              muxOutConnector[16] = fifoOut[3][8];
              muxOutConnector[17] = fifoOut[4][8];
              muxOutConnector[18] = fifoOut[5][8];
              muxOutConnector[19] = fifoOut[6][8];
              muxOutConnector[20] = fifoOut[7][8];
              muxOutConnector[21] = fifoOut[8][8];
              muxOutConnector[22] = fifoOut[9][8];
              muxOutConnector[23] = fifoOut[10][8];
              muxOutConnector[24] = fifoOut[11][8];
              muxOutConnector[25] = fifoOut[12][8];
              muxOutConnector[26] = fifoOut[45][2];
              muxOutConnector[27] = fifoOut[46][2];
              muxOutConnector[28] = fifoOut[47][2];
              muxOutConnector[29] = fifoOut[48][2];
              muxOutConnector[30] = fifoOut[49][2];
              muxOutConnector[31] = fifoOut[50][2];
              muxOutConnector[32] = fifoOut[51][2];
              muxOutConnector[33] = fifoOut[26][1];
              muxOutConnector[34] = fifoOut[27][1];
              muxOutConnector[35] = fifoOut[28][1];
              muxOutConnector[36] = fifoOut[29][1];
              muxOutConnector[37] = fifoOut[30][1];
              muxOutConnector[38] = fifoOut[31][1];
              muxOutConnector[39] = fifoOut[32][1];
              muxOutConnector[40] = fifoOut[33][1];
              muxOutConnector[41] = fifoOut[34][1];
              muxOutConnector[42] = fifoOut[35][1];
              muxOutConnector[43] = fifoOut[36][1];
              muxOutConnector[44] = fifoOut[37][1];
              muxOutConnector[45] = fifoOut[38][1];
              muxOutConnector[46] = fifoOut[39][1];
              muxOutConnector[47] = fifoOut[40][1];
              muxOutConnector[48] = fifoOut[41][1];
              muxOutConnector[49] = fifoOut[42][1];
              muxOutConnector[50] = fifoOut[43][1];
              muxOutConnector[51] = fifoOut[44][1];
       end
       7: begin
              muxOutConnector[0] = fifoOut[13][9];
              muxOutConnector[1] = fifoOut[14][9];
              muxOutConnector[2] = fifoOut[15][9];
              muxOutConnector[3] = fifoOut[16][9];
              muxOutConnector[4] = fifoOut[17][9];
              muxOutConnector[5] = fifoOut[18][9];
              muxOutConnector[6] = fifoOut[19][9];
              muxOutConnector[7] = fifoOut[20][9];
              muxOutConnector[8] = fifoOut[21][9];
              muxOutConnector[9] = fifoOut[22][9];
              muxOutConnector[10] = fifoOut[23][9];
              muxOutConnector[11] = fifoOut[24][9];
              muxOutConnector[12] = fifoOut[25][9];
              muxOutConnector[13] = fifoOut[0][8];
              muxOutConnector[14] = fifoOut[1][8];
              muxOutConnector[15] = fifoOut[2][8];
              muxOutConnector[16] = fifoOut[3][8];
              muxOutConnector[17] = fifoOut[4][8];
              muxOutConnector[18] = fifoOut[5][8];
              muxOutConnector[19] = fifoOut[6][8];
              muxOutConnector[20] = fifoOut[7][8];
              muxOutConnector[21] = fifoOut[8][8];
              muxOutConnector[22] = fifoOut[9][8];
              muxOutConnector[23] = fifoOut[10][8];
              muxOutConnector[24] = fifoOut[11][8];
              muxOutConnector[25] = fifoOut[12][8];
              muxOutConnector[26] = fifoOut[45][2];
              muxOutConnector[27] = fifoOut[46][2];
              muxOutConnector[28] = fifoOut[47][2];
              muxOutConnector[29] = fifoOut[48][2];
              muxOutConnector[30] = fifoOut[49][2];
              muxOutConnector[31] = fifoOut[50][2];
              muxOutConnector[32] = fifoOut[51][2];
              muxOutConnector[33] = fifoOut[26][1];
              muxOutConnector[34] = fifoOut[27][1];
              muxOutConnector[35] = fifoOut[28][1];
              muxOutConnector[36] = fifoOut[29][1];
              muxOutConnector[37] = fifoOut[30][1];
              muxOutConnector[38] = fifoOut[31][1];
              muxOutConnector[39] = fifoOut[32][1];
              muxOutConnector[40] = fifoOut[33][1];
              muxOutConnector[41] = fifoOut[34][1];
              muxOutConnector[42] = fifoOut[35][1];
              muxOutConnector[43] = fifoOut[36][1];
              muxOutConnector[44] = fifoOut[37][1];
              muxOutConnector[45] = fifoOut[38][1];
              muxOutConnector[46] = fifoOut[39][1];
              muxOutConnector[47] = fifoOut[40][1];
              muxOutConnector[48] = fifoOut[41][1];
              muxOutConnector[49] = fifoOut[42][1];
              muxOutConnector[50] = fifoOut[43][1];
              muxOutConnector[51] = fifoOut[44][1];
       end
       8: begin
              muxOutConnector[0] = fifoOut[13][9];
              muxOutConnector[1] = fifoOut[14][9];
              muxOutConnector[2] = fifoOut[15][9];
              muxOutConnector[3] = fifoOut[16][9];
              muxOutConnector[4] = fifoOut[17][9];
              muxOutConnector[5] = fifoOut[18][9];
              muxOutConnector[6] = fifoOut[19][9];
              muxOutConnector[7] = fifoOut[20][9];
              muxOutConnector[8] = fifoOut[21][9];
              muxOutConnector[9] = fifoOut[22][9];
              muxOutConnector[10] = fifoOut[23][9];
              muxOutConnector[11] = fifoOut[24][9];
              muxOutConnector[12] = fifoOut[25][9];
              muxOutConnector[13] = fifoOut[0][8];
              muxOutConnector[14] = fifoOut[1][8];
              muxOutConnector[15] = fifoOut[2][8];
              muxOutConnector[16] = fifoOut[3][8];
              muxOutConnector[17] = fifoOut[4][8];
              muxOutConnector[18] = fifoOut[5][8];
              muxOutConnector[19] = fifoOut[6][8];
              muxOutConnector[20] = fifoOut[7][8];
              muxOutConnector[21] = fifoOut[8][8];
              muxOutConnector[22] = fifoOut[9][8];
              muxOutConnector[23] = fifoOut[10][8];
              muxOutConnector[24] = fifoOut[11][8];
              muxOutConnector[25] = fifoOut[12][8];
              muxOutConnector[26] = fifoOut[45][2];
              muxOutConnector[27] = fifoOut[46][2];
              muxOutConnector[28] = fifoOut[47][2];
              muxOutConnector[29] = fifoOut[48][2];
              muxOutConnector[30] = fifoOut[49][2];
              muxOutConnector[31] = fifoOut[50][2];
              muxOutConnector[32] = fifoOut[51][2];
              muxOutConnector[33] = fifoOut[26][1];
              muxOutConnector[34] = fifoOut[27][1];
              muxOutConnector[35] = fifoOut[28][1];
              muxOutConnector[36] = fifoOut[29][1];
              muxOutConnector[37] = fifoOut[30][1];
              muxOutConnector[38] = fifoOut[31][1];
              muxOutConnector[39] = fifoOut[32][1];
              muxOutConnector[40] = fifoOut[33][1];
              muxOutConnector[41] = fifoOut[34][1];
              muxOutConnector[42] = fifoOut[35][1];
              muxOutConnector[43] = fifoOut[36][1];
              muxOutConnector[44] = fifoOut[37][1];
              muxOutConnector[45] = fifoOut[38][1];
              muxOutConnector[46] = fifoOut[39][1];
              muxOutConnector[47] = fifoOut[40][1];
              muxOutConnector[48] = fifoOut[41][1];
              muxOutConnector[49] = fifoOut[42][1];
              muxOutConnector[50] = fifoOut[43][1];
              muxOutConnector[51] = fifoOut[44][1];
       end
       9: begin
              muxOutConnector[0] = fifoOut[13][9];
              muxOutConnector[1] = fifoOut[14][9];
              muxOutConnector[2] = fifoOut[15][9];
              muxOutConnector[3] = fifoOut[16][9];
              muxOutConnector[4] = fifoOut[48][8];
              muxOutConnector[5] = fifoOut[49][8];
              muxOutConnector[6] = fifoOut[50][8];
              muxOutConnector[7] = fifoOut[51][8];
              muxOutConnector[8] = fifoOut[26][7];
              muxOutConnector[9] = fifoOut[27][7];
              muxOutConnector[10] = fifoOut[28][7];
              muxOutConnector[11] = fifoOut[29][7];
              muxOutConnector[12] = fifoOut[30][7];
              muxOutConnector[13] = fifoOut[31][7];
              muxOutConnector[14] = fifoOut[32][7];
              muxOutConnector[15] = fifoOut[33][7];
              muxOutConnector[16] = fifoOut[34][7];
              muxOutConnector[17] = fifoOut[35][7];
              muxOutConnector[18] = fifoOut[36][7];
              muxOutConnector[19] = fifoOut[37][7];
              muxOutConnector[20] = fifoOut[38][7];
              muxOutConnector[21] = fifoOut[39][7];
              muxOutConnector[22] = fifoOut[40][7];
              muxOutConnector[23] = fifoOut[41][7];
              muxOutConnector[24] = fifoOut[42][7];
              muxOutConnector[25] = fifoOut[43][7];
              muxOutConnector[26] = fifoOut[45][2];
              muxOutConnector[27] = fifoOut[46][2];
              muxOutConnector[28] = fifoOut[47][2];
              muxOutConnector[29] = fifoOut[48][2];
              muxOutConnector[30] = fifoOut[49][2];
              muxOutConnector[31] = fifoOut[50][2];
              muxOutConnector[32] = fifoOut[51][2];
              muxOutConnector[33] = fifoOut[26][1];
              muxOutConnector[34] = fifoOut[27][1];
              muxOutConnector[35] = fifoOut[28][1];
              muxOutConnector[36] = fifoOut[29][1];
              muxOutConnector[37] = fifoOut[30][1];
              muxOutConnector[38] = fifoOut[31][1];
              muxOutConnector[39] = fifoOut[32][1];
              muxOutConnector[40] = fifoOut[33][1];
              muxOutConnector[41] = fifoOut[34][1];
              muxOutConnector[42] = fifoOut[35][1];
              muxOutConnector[43] = fifoOut[36][1];
              muxOutConnector[44] = fifoOut[37][1];
              muxOutConnector[45] = fifoOut[38][1];
              muxOutConnector[46] = fifoOut[39][1];
              muxOutConnector[47] = fifoOut[40][1];
              muxOutConnector[48] = fifoOut[41][1];
              muxOutConnector[49] = fifoOut[42][1];
              muxOutConnector[50] = fifoOut[43][1];
              muxOutConnector[51] = fifoOut[44][1];
       end
       10: begin
              muxOutConnector[0] = fifoOut[44][8];
              muxOutConnector[1] = fifoOut[45][8];
              muxOutConnector[2] = fifoOut[46][8];
              muxOutConnector[3] = fifoOut[47][8];
              muxOutConnector[4] = fifoOut[48][8];
              muxOutConnector[5] = fifoOut[49][8];
              muxOutConnector[6] = fifoOut[50][8];
              muxOutConnector[7] = fifoOut[51][8];
              muxOutConnector[8] = fifoOut[26][7];
              muxOutConnector[9] = fifoOut[27][7];
              muxOutConnector[10] = fifoOut[28][7];
              muxOutConnector[11] = fifoOut[29][7];
              muxOutConnector[12] = fifoOut[30][7];
              muxOutConnector[13] = fifoOut[31][7];
              muxOutConnector[14] = fifoOut[32][7];
              muxOutConnector[15] = fifoOut[33][7];
              muxOutConnector[16] = fifoOut[34][7];
              muxOutConnector[17] = fifoOut[35][7];
              muxOutConnector[18] = fifoOut[36][7];
              muxOutConnector[19] = fifoOut[37][7];
              muxOutConnector[20] = fifoOut[38][7];
              muxOutConnector[21] = fifoOut[39][7];
              muxOutConnector[22] = fifoOut[40][7];
              muxOutConnector[23] = fifoOut[41][7];
              muxOutConnector[24] = fifoOut[42][7];
              muxOutConnector[25] = fifoOut[43][7];
              muxOutConnector[26] = fifoOut[45][2];
              muxOutConnector[27] = fifoOut[46][2];
              muxOutConnector[28] = fifoOut[47][2];
              muxOutConnector[29] = fifoOut[0][9];
              muxOutConnector[30] = fifoOut[1][9];
              muxOutConnector[31] = fifoOut[2][9];
              muxOutConnector[32] = fifoOut[3][9];
              muxOutConnector[33] = fifoOut[4][9];
              muxOutConnector[34] = fifoOut[5][9];
              muxOutConnector[35] = fifoOut[6][9];
              muxOutConnector[36] = fifoOut[7][9];
              muxOutConnector[37] = fifoOut[8][9];
              muxOutConnector[38] = fifoOut[9][9];
              muxOutConnector[39] = fifoOut[10][9];
              muxOutConnector[40] = fifoOut[11][9];
              muxOutConnector[41] = fifoOut[12][9];
              muxOutConnector[42] = fifoOut[13][9];
              muxOutConnector[43] = fifoOut[14][9];
              muxOutConnector[44] = fifoOut[15][9];
              muxOutConnector[45] = fifoOut[16][9];
              muxOutConnector[46] = fifoOut[17][9];
              muxOutConnector[47] = fifoOut[18][9];
              muxOutConnector[48] = fifoOut[19][9];
              muxOutConnector[49] = fifoOut[20][9];
              muxOutConnector[50] = fifoOut[21][9];
              muxOutConnector[51] = fifoOut[22][9];
       end
       11: begin
              muxOutConnector[0] = fifoOut[44][8];
              muxOutConnector[1] = fifoOut[45][8];
              muxOutConnector[2] = fifoOut[46][8];
              muxOutConnector[3] = fifoOut[47][8];
              muxOutConnector[4] = fifoOut[48][8];
              muxOutConnector[5] = fifoOut[49][8];
              muxOutConnector[6] = fifoOut[50][8];
              muxOutConnector[7] = fifoOut[51][8];
              muxOutConnector[8] = fifoOut[26][7];
              muxOutConnector[9] = fifoOut[27][7];
              muxOutConnector[10] = fifoOut[28][7];
              muxOutConnector[11] = fifoOut[29][7];
              muxOutConnector[12] = fifoOut[30][7];
              muxOutConnector[13] = fifoOut[31][7];
              muxOutConnector[14] = fifoOut[32][7];
              muxOutConnector[15] = fifoOut[33][7];
              muxOutConnector[16] = fifoOut[34][7];
              muxOutConnector[17] = fifoOut[35][7];
              muxOutConnector[18] = fifoOut[36][7];
              muxOutConnector[19] = fifoOut[37][7];
              muxOutConnector[20] = fifoOut[38][7];
              muxOutConnector[21] = fifoOut[39][7];
              muxOutConnector[22] = fifoOut[40][7];
              muxOutConnector[23] = fifoOut[41][7];
              muxOutConnector[24] = fifoOut[42][7];
              muxOutConnector[25] = fifoOut[43][7];
              muxOutConnector[26] = fifoOut[23][10];
              muxOutConnector[27] = fifoOut[24][10];
              muxOutConnector[28] = fifoOut[25][10];
              muxOutConnector[29] = fifoOut[0][9];
              muxOutConnector[30] = fifoOut[1][9];
              muxOutConnector[31] = fifoOut[2][9];
              muxOutConnector[32] = fifoOut[3][9];
              muxOutConnector[33] = fifoOut[4][9];
              muxOutConnector[34] = fifoOut[5][9];
              muxOutConnector[35] = fifoOut[6][9];
              muxOutConnector[36] = fifoOut[7][9];
              muxOutConnector[37] = fifoOut[8][9];
              muxOutConnector[38] = fifoOut[9][9];
              muxOutConnector[39] = fifoOut[10][9];
              muxOutConnector[40] = fifoOut[11][9];
              muxOutConnector[41] = fifoOut[12][9];
              muxOutConnector[42] = fifoOut[13][9];
              muxOutConnector[43] = fifoOut[14][9];
              muxOutConnector[44] = fifoOut[15][9];
              muxOutConnector[45] = fifoOut[16][9];
              muxOutConnector[46] = fifoOut[17][9];
              muxOutConnector[47] = fifoOut[18][9];
              muxOutConnector[48] = fifoOut[19][9];
              muxOutConnector[49] = fifoOut[20][9];
              muxOutConnector[50] = fifoOut[21][9];
              muxOutConnector[51] = fifoOut[22][9];
       end
       12: begin
              muxOutConnector[0] = fifoOut[44][8];
              muxOutConnector[1] = fifoOut[45][8];
              muxOutConnector[2] = fifoOut[46][8];
              muxOutConnector[3] = fifoOut[47][8];
              muxOutConnector[4] = fifoOut[48][8];
              muxOutConnector[5] = fifoOut[49][8];
              muxOutConnector[6] = fifoOut[50][8];
              muxOutConnector[7] = fifoOut[51][8];
              muxOutConnector[8] = fifoOut[26][7];
              muxOutConnector[9] = fifoOut[27][7];
              muxOutConnector[10] = fifoOut[28][7];
              muxOutConnector[11] = fifoOut[29][7];
              muxOutConnector[12] = fifoOut[30][7];
              muxOutConnector[13] = fifoOut[31][7];
              muxOutConnector[14] = fifoOut[32][7];
              muxOutConnector[15] = fifoOut[33][7];
              muxOutConnector[16] = fifoOut[34][7];
              muxOutConnector[17] = fifoOut[35][7];
              muxOutConnector[18] = fifoOut[36][7];
              muxOutConnector[19] = fifoOut[37][7];
              muxOutConnector[20] = fifoOut[38][7];
              muxOutConnector[21] = fifoOut[39][7];
              muxOutConnector[22] = fifoOut[40][7];
              muxOutConnector[23] = fifoOut[41][7];
              muxOutConnector[24] = fifoOut[42][7];
              muxOutConnector[25] = fifoOut[43][7];
              muxOutConnector[26] = fifoOut[23][10];
              muxOutConnector[27] = fifoOut[24][10];
              muxOutConnector[28] = fifoOut[25][10];
              muxOutConnector[29] = fifoOut[0][9];
              muxOutConnector[30] = fifoOut[1][9];
              muxOutConnector[31] = fifoOut[2][9];
              muxOutConnector[32] = fifoOut[3][9];
              muxOutConnector[33] = fifoOut[4][9];
              muxOutConnector[34] = fifoOut[5][9];
              muxOutConnector[35] = fifoOut[6][9];
              muxOutConnector[36] = fifoOut[7][9];
              muxOutConnector[37] = fifoOut[8][9];
              muxOutConnector[38] = fifoOut[9][9];
              muxOutConnector[39] = fifoOut[10][9];
              muxOutConnector[40] = fifoOut[11][9];
              muxOutConnector[41] = fifoOut[12][9];
              muxOutConnector[42] = fifoOut[13][9];
              muxOutConnector[43] = fifoOut[14][9];
              muxOutConnector[44] = fifoOut[15][9];
              muxOutConnector[45] = fifoOut[16][9];
              muxOutConnector[46] = fifoOut[17][9];
              muxOutConnector[47] = fifoOut[18][9];
              muxOutConnector[48] = fifoOut[19][9];
              muxOutConnector[49] = fifoOut[20][9];
              muxOutConnector[50] = fifoOut[21][9];
              muxOutConnector[51] = fifoOut[22][9];
       end
       13: begin
              muxOutConnector[0] = fifoOut[44][8];
              muxOutConnector[1] = fifoOut[45][8];
              muxOutConnector[2] = fifoOut[46][8];
              muxOutConnector[3] = fifoOut[47][8];
              muxOutConnector[4] = fifoOut[48][8];
              muxOutConnector[5] = fifoOut[49][8];
              muxOutConnector[6] = fifoOut[50][8];
              muxOutConnector[7] = fifoOut[51][8];
              muxOutConnector[8] = fifoOut[26][7];
              muxOutConnector[9] = fifoOut[27][7];
              muxOutConnector[10] = fifoOut[28][7];
              muxOutConnector[11] = fifoOut[29][7];
              muxOutConnector[12] = fifoOut[30][7];
              muxOutConnector[13] = fifoOut[31][7];
              muxOutConnector[14] = fifoOut[32][7];
              muxOutConnector[15] = fifoOut[33][7];
              muxOutConnector[16] = fifoOut[34][7];
              muxOutConnector[17] = fifoOut[35][7];
              muxOutConnector[18] = fifoOut[36][7];
              muxOutConnector[19] = fifoOut[37][7];
              muxOutConnector[20] = fifoOut[38][7];
              muxOutConnector[21] = fifoOut[39][7];
              muxOutConnector[22] = fifoOut[40][7];
              muxOutConnector[23] = fifoOut[41][7];
              muxOutConnector[24] = fifoOut[42][7];
              muxOutConnector[25] = fifoOut[43][7];
              muxOutConnector[26] = fifoOut[23][10];
              muxOutConnector[27] = fifoOut[24][10];
              muxOutConnector[28] = fifoOut[25][10];
              muxOutConnector[29] = fifoOut[0][9];
              muxOutConnector[30] = fifoOut[1][9];
              muxOutConnector[31] = fifoOut[2][9];
              muxOutConnector[32] = fifoOut[3][9];
              muxOutConnector[33] = fifoOut[4][9];
              muxOutConnector[34] = fifoOut[5][9];
              muxOutConnector[35] = fifoOut[6][9];
              muxOutConnector[36] = fifoOut[7][9];
              muxOutConnector[37] = fifoOut[8][9];
              muxOutConnector[38] = fifoOut[9][9];
              muxOutConnector[39] = fifoOut[10][9];
              muxOutConnector[40] = fifoOut[11][9];
              muxOutConnector[41] = fifoOut[12][9];
              muxOutConnector[42] = fifoOut[13][9];
              muxOutConnector[43] = fifoOut[14][9];
              muxOutConnector[44] = fifoOut[15][9];
              muxOutConnector[45] = fifoOut[16][9];
              muxOutConnector[46] = fifoOut[17][9];
              muxOutConnector[47] = fifoOut[18][9];
              muxOutConnector[48] = fifoOut[19][9];
              muxOutConnector[49] = fifoOut[20][9];
              muxOutConnector[50] = fifoOut[21][9];
              muxOutConnector[51] = fifoOut[22][9];
       end
       14: begin
              muxOutConnector[0] = fifoOut[44][8];
              muxOutConnector[1] = fifoOut[45][8];
              muxOutConnector[2] = fifoOut[46][8];
              muxOutConnector[3] = fifoOut[47][8];
              muxOutConnector[4] = fifoOut[48][8];
              muxOutConnector[5] = fifoOut[49][8];
              muxOutConnector[6] = fifoOut[50][8];
              muxOutConnector[7] = fifoOut[51][8];
              muxOutConnector[8] = fifoOut[26][7];
              muxOutConnector[9] = fifoOut[27][7];
              muxOutConnector[10] = fifoOut[28][7];
              muxOutConnector[11] = fifoOut[29][7];
              muxOutConnector[12] = fifoOut[30][7];
              muxOutConnector[13] = fifoOut[31][7];
              muxOutConnector[14] = fifoOut[32][7];
              muxOutConnector[15] = fifoOut[33][7];
              muxOutConnector[16] = fifoOut[34][7];
              muxOutConnector[17] = fifoOut[35][7];
              muxOutConnector[18] = fifoOut[36][7];
              muxOutConnector[19] = fifoOut[37][7];
              muxOutConnector[20] = fifoOut[38][7];
              muxOutConnector[21] = fifoOut[39][7];
              muxOutConnector[22] = fifoOut[40][7];
              muxOutConnector[23] = fifoOut[41][7];
              muxOutConnector[24] = fifoOut[42][7];
              muxOutConnector[25] = fifoOut[43][7];
              muxOutConnector[26] = fifoOut[23][10];
              muxOutConnector[27] = fifoOut[24][10];
              muxOutConnector[28] = fifoOut[25][10];
              muxOutConnector[29] = fifoOut[0][9];
              muxOutConnector[30] = fifoOut[1][9];
              muxOutConnector[31] = fifoOut[2][9];
              muxOutConnector[32] = fifoOut[3][9];
              muxOutConnector[33] = fifoOut[4][9];
              muxOutConnector[34] = fifoOut[5][9];
              muxOutConnector[35] = fifoOut[6][9];
              muxOutConnector[36] = fifoOut[7][9];
              muxOutConnector[37] = fifoOut[8][9];
              muxOutConnector[38] = fifoOut[9][9];
              muxOutConnector[39] = fifoOut[10][9];
              muxOutConnector[40] = fifoOut[11][9];
              muxOutConnector[41] = fifoOut[12][9];
              muxOutConnector[42] = fifoOut[13][9];
              muxOutConnector[43] = fifoOut[14][9];
              muxOutConnector[44] = fifoOut[15][9];
              muxOutConnector[45] = fifoOut[16][9];
              muxOutConnector[46] = fifoOut[17][9];
              muxOutConnector[47] = fifoOut[18][9];
              muxOutConnector[48] = fifoOut[19][9];
              muxOutConnector[49] = fifoOut[20][9];
              muxOutConnector[50] = fifoOut[21][9];
              muxOutConnector[51] = fifoOut[22][9];
       end
       15: begin
              muxOutConnector[0] = fifoOut[44][8];
              muxOutConnector[1] = fifoOut[45][8];
              muxOutConnector[2] = fifoOut[46][8];
              muxOutConnector[3] = fifoOut[47][8];
              muxOutConnector[4] = fifoOut[48][8];
              muxOutConnector[5] = fifoOut[49][8];
              muxOutConnector[6] = fifoOut[50][8];
              muxOutConnector[7] = fifoOut[51][8];
              muxOutConnector[8] = fifoOut[26][7];
              muxOutConnector[9] = fifoOut[27][7];
              muxOutConnector[10] = fifoOut[28][7];
              muxOutConnector[11] = fifoOut[29][7];
              muxOutConnector[12] = fifoOut[30][7];
              muxOutConnector[13] = fifoOut[31][7];
              muxOutConnector[14] = fifoOut[32][7];
              muxOutConnector[15] = fifoOut[33][7];
              muxOutConnector[16] = fifoOut[34][7];
              muxOutConnector[17] = fifoOut[35][7];
              muxOutConnector[18] = fifoOut[36][7];
              muxOutConnector[19] = fifoOut[37][7];
              muxOutConnector[20] = fifoOut[38][7];
              muxOutConnector[21] = fifoOut[39][7];
              muxOutConnector[22] = fifoOut[40][7];
              muxOutConnector[23] = fifoOut[41][7];
              muxOutConnector[24] = fifoOut[42][7];
              muxOutConnector[25] = fifoOut[43][7];
              muxOutConnector[26] = fifoOut[23][10];
              muxOutConnector[27] = fifoOut[24][10];
              muxOutConnector[28] = fifoOut[25][10];
              muxOutConnector[29] = fifoOut[0][9];
              muxOutConnector[30] = fifoOut[1][9];
              muxOutConnector[31] = fifoOut[2][9];
              muxOutConnector[32] = fifoOut[3][9];
              muxOutConnector[33] = fifoOut[4][9];
              muxOutConnector[34] = fifoOut[5][9];
              muxOutConnector[35] = fifoOut[6][9];
              muxOutConnector[36] = fifoOut[7][9];
              muxOutConnector[37] = fifoOut[8][9];
              muxOutConnector[38] = fifoOut[9][9];
              muxOutConnector[39] = fifoOut[10][9];
              muxOutConnector[40] = fifoOut[11][9];
              muxOutConnector[41] = fifoOut[12][9];
              muxOutConnector[42] = fifoOut[13][9];
              muxOutConnector[43] = fifoOut[14][9];
              muxOutConnector[44] = fifoOut[15][9];
              muxOutConnector[45] = fifoOut[16][9];
              muxOutConnector[46] = fifoOut[17][9];
              muxOutConnector[47] = fifoOut[18][9];
              muxOutConnector[48] = fifoOut[19][9];
              muxOutConnector[49] = fifoOut[20][9];
              muxOutConnector[50] = fifoOut[21][9];
              muxOutConnector[51] = fifoOut[22][9];
       end
       16: begin
              muxOutConnector[0] = fifoOut[44][8];
              muxOutConnector[1] = fifoOut[45][8];
              muxOutConnector[2] = fifoOut[46][8];
              muxOutConnector[3] = fifoOut[47][8];
              muxOutConnector[4] = fifoOut[48][8];
              muxOutConnector[5] = fifoOut[49][8];
              muxOutConnector[6] = fifoOut[50][8];
              muxOutConnector[7] = fifoOut[51][8];
              muxOutConnector[8] = fifoOut[26][7];
              muxOutConnector[9] = fifoOut[27][7];
              muxOutConnector[10] = fifoOut[28][7];
              muxOutConnector[11] = fifoOut[29][7];
              muxOutConnector[12] = fifoOut[30][7];
              muxOutConnector[13] = fifoOut[31][7];
              muxOutConnector[14] = fifoOut[32][7];
              muxOutConnector[15] = fifoOut[33][7];
              muxOutConnector[16] = fifoOut[34][7];
              muxOutConnector[17] = fifoOut[35][7];
              muxOutConnector[18] = fifoOut[36][7];
              muxOutConnector[19] = fifoOut[37][7];
              muxOutConnector[20] = fifoOut[38][7];
              muxOutConnector[21] = fifoOut[39][7];
              muxOutConnector[22] = fifoOut[40][7];
              muxOutConnector[23] = fifoOut[41][7];
              muxOutConnector[24] = fifoOut[42][7];
              muxOutConnector[25] = fifoOut[43][7];
              muxOutConnector[26] = fifoOut[23][10];
              muxOutConnector[27] = fifoOut[24][10];
              muxOutConnector[28] = fifoOut[25][10];
              muxOutConnector[29] = fifoOut[0][9];
              muxOutConnector[30] = fifoOut[1][9];
              muxOutConnector[31] = fifoOut[2][9];
              muxOutConnector[32] = fifoOut[3][9];
              muxOutConnector[33] = fifoOut[4][9];
              muxOutConnector[34] = fifoOut[5][9];
              muxOutConnector[35] = fifoOut[6][9];
              muxOutConnector[36] = fifoOut[7][9];
              muxOutConnector[37] = fifoOut[8][9];
              muxOutConnector[38] = fifoOut[9][9];
              muxOutConnector[39] = fifoOut[10][9];
              muxOutConnector[40] = fifoOut[11][9];
              muxOutConnector[41] = fifoOut[12][9];
              muxOutConnector[42] = fifoOut[13][9];
              muxOutConnector[43] = fifoOut[14][9];
              muxOutConnector[44] = fifoOut[15][9];
              muxOutConnector[45] = fifoOut[16][9];
              muxOutConnector[46] = fifoOut[17][9];
              muxOutConnector[47] = fifoOut[18][9];
              muxOutConnector[48] = fifoOut[19][9];
              muxOutConnector[49] = fifoOut[20][9];
              muxOutConnector[50] = fifoOut[21][9];
              muxOutConnector[51] = fifoOut[22][9];
       end
       17: begin
              muxOutConnector[0] = fifoOut[44][8];
              muxOutConnector[1] = fifoOut[45][8];
              muxOutConnector[2] = fifoOut[46][8];
              muxOutConnector[3] = fifoOut[47][8];
              muxOutConnector[4] = fifoOut[48][8];
              muxOutConnector[5] = fifoOut[49][8];
              muxOutConnector[6] = fifoOut[50][8];
              muxOutConnector[7] = fifoOut[51][8];
              muxOutConnector[8] = fifoOut[26][7];
              muxOutConnector[9] = fifoOut[27][7];
              muxOutConnector[10] = fifoOut[28][7];
              muxOutConnector[11] = fifoOut[29][7];
              muxOutConnector[12] = fifoOut[30][7];
              muxOutConnector[13] = fifoOut[31][7];
              muxOutConnector[14] = fifoOut[32][7];
              muxOutConnector[15] = fifoOut[33][7];
              muxOutConnector[16] = fifoOut[34][7];
              muxOutConnector[17] = fifoOut[35][7];
              muxOutConnector[18] = fifoOut[36][7];
              muxOutConnector[19] = fifoOut[37][7];
              muxOutConnector[20] = fifoOut[38][7];
              muxOutConnector[21] = fifoOut[39][7];
              muxOutConnector[22] = fifoOut[40][7];
              muxOutConnector[23] = fifoOut[41][7];
              muxOutConnector[24] = fifoOut[42][7];
              muxOutConnector[25] = fifoOut[43][7];
              muxOutConnector[26] = fifoOut[23][10];
              muxOutConnector[27] = fifoOut[24][10];
              muxOutConnector[28] = fifoOut[25][10];
              muxOutConnector[29] = fifoOut[0][9];
              muxOutConnector[30] = fifoOut[1][9];
              muxOutConnector[31] = fifoOut[2][9];
              muxOutConnector[32] = fifoOut[3][9];
              muxOutConnector[33] = fifoOut[4][9];
              muxOutConnector[34] = fifoOut[5][9];
              muxOutConnector[35] = fifoOut[6][9];
              muxOutConnector[36] = fifoOut[7][9];
              muxOutConnector[37] = fifoOut[8][9];
              muxOutConnector[38] = fifoOut[9][9];
              muxOutConnector[39] = fifoOut[10][9];
              muxOutConnector[40] = fifoOut[11][9];
              muxOutConnector[41] = fifoOut[12][9];
              muxOutConnector[42] = fifoOut[13][9];
              muxOutConnector[43] = fifoOut[14][9];
              muxOutConnector[44] = fifoOut[15][9];
              muxOutConnector[45] = fifoOut[16][9];
              muxOutConnector[46] = fifoOut[17][9];
              muxOutConnector[47] = fifoOut[18][9];
              muxOutConnector[48] = fifoOut[19][9];
              muxOutConnector[49] = fifoOut[20][9];
              muxOutConnector[50] = fifoOut[21][9];
              muxOutConnector[51] = fifoOut[22][9];
       end
       18: begin
              muxOutConnector[0] = fifoOut[44][8];
              muxOutConnector[1] = fifoOut[45][8];
              muxOutConnector[2] = fifoOut[46][8];
              muxOutConnector[3] = fifoOut[47][8];
              muxOutConnector[4] = fifoOut[48][8];
              muxOutConnector[5] = fifoOut[49][8];
              muxOutConnector[6] = fifoOut[50][8];
              muxOutConnector[7] = fifoOut[51][8];
              muxOutConnector[8] = fifoOut[26][7];
              muxOutConnector[9] = fifoOut[27][7];
              muxOutConnector[10] = fifoOut[28][7];
              muxOutConnector[11] = fifoOut[29][7];
              muxOutConnector[12] = fifoOut[30][7];
              muxOutConnector[13] = fifoOut[31][7];
              muxOutConnector[14] = fifoOut[32][7];
              muxOutConnector[15] = fifoOut[33][7];
              muxOutConnector[16] = fifoOut[34][7];
              muxOutConnector[17] = fifoOut[35][7];
              muxOutConnector[18] = fifoOut[36][7];
              muxOutConnector[19] = fifoOut[37][7];
              muxOutConnector[20] = fifoOut[38][7];
              muxOutConnector[21] = fifoOut[39][7];
              muxOutConnector[22] = fifoOut[40][7];
              muxOutConnector[23] = fifoOut[41][7];
              muxOutConnector[24] = fifoOut[42][7];
              muxOutConnector[25] = fifoOut[43][7];
              muxOutConnector[26] = fifoOut[23][10];
              muxOutConnector[27] = fifoOut[24][10];
              muxOutConnector[28] = fifoOut[25][10];
              muxOutConnector[29] = fifoOut[0][9];
              muxOutConnector[30] = fifoOut[1][9];
              muxOutConnector[31] = fifoOut[2][9];
              muxOutConnector[32] = fifoOut[3][9];
              muxOutConnector[33] = fifoOut[4][9];
              muxOutConnector[34] = fifoOut[5][9];
              muxOutConnector[35] = fifoOut[6][9];
              muxOutConnector[36] = fifoOut[7][9];
              muxOutConnector[37] = fifoOut[8][9];
              muxOutConnector[38] = fifoOut[9][9];
              muxOutConnector[39] = fifoOut[10][9];
              muxOutConnector[40] = fifoOut[11][9];
              muxOutConnector[41] = fifoOut[12][9];
              muxOutConnector[42] = fifoOut[13][9];
              muxOutConnector[43] = fifoOut[14][9];
              muxOutConnector[44] = fifoOut[15][9];
              muxOutConnector[45] = fifoOut[16][9];
              muxOutConnector[46] = fifoOut[17][9];
              muxOutConnector[47] = fifoOut[18][9];
              muxOutConnector[48] = fifoOut[19][9];
              muxOutConnector[49] = fifoOut[20][9];
              muxOutConnector[50] = fifoOut[21][9];
              muxOutConnector[51] = fifoOut[22][9];
       end
       19: begin
              muxOutConnector[0] = fifoOut[44][8];
              muxOutConnector[1] = fifoOut[45][8];
              muxOutConnector[2] = fifoOut[46][8];
              muxOutConnector[3] = fifoOut[47][8];
              muxOutConnector[4] = fifoOut[48][8];
              muxOutConnector[5] = fifoOut[49][8];
              muxOutConnector[6] = fifoOut[50][8];
              muxOutConnector[7] = fifoOut[51][8];
              muxOutConnector[8] = fifoOut[26][7];
              muxOutConnector[9] = fifoOut[27][7];
              muxOutConnector[10] = fifoOut[28][7];
              muxOutConnector[11] = fifoOut[29][7];
              muxOutConnector[12] = fifoOut[30][7];
              muxOutConnector[13] = fifoOut[31][7];
              muxOutConnector[14] = fifoOut[32][7];
              muxOutConnector[15] = fifoOut[33][7];
              muxOutConnector[16] = fifoOut[34][7];
              muxOutConnector[17] = maxVal;
              muxOutConnector[18] = maxVal;
              muxOutConnector[19] = maxVal;
              muxOutConnector[20] = maxVal;
              muxOutConnector[21] = maxVal;
              muxOutConnector[22] = maxVal;
              muxOutConnector[23] = maxVal;
              muxOutConnector[24] = maxVal;
              muxOutConnector[25] = maxVal;
              muxOutConnector[26] = fifoOut[23][10];
              muxOutConnector[27] = fifoOut[24][10];
              muxOutConnector[28] = fifoOut[25][10];
              muxOutConnector[29] = fifoOut[0][9];
              muxOutConnector[30] = fifoOut[1][9];
              muxOutConnector[31] = fifoOut[2][9];
              muxOutConnector[32] = fifoOut[3][9];
              muxOutConnector[33] = fifoOut[4][9];
              muxOutConnector[34] = fifoOut[5][9];
              muxOutConnector[35] = fifoOut[6][9];
              muxOutConnector[36] = fifoOut[7][9];
              muxOutConnector[37] = fifoOut[8][9];
              muxOutConnector[38] = fifoOut[9][9];
              muxOutConnector[39] = fifoOut[10][9];
              muxOutConnector[40] = fifoOut[11][9];
              muxOutConnector[41] = fifoOut[12][9];
              muxOutConnector[42] = fifoOut[13][9];
              muxOutConnector[43] = maxVal;
              muxOutConnector[44] = maxVal;
              muxOutConnector[45] = maxVal;
              muxOutConnector[46] = maxVal;
              muxOutConnector[47] = maxVal;
              muxOutConnector[48] = maxVal;
              muxOutConnector[49] = maxVal;
              muxOutConnector[50] = maxVal;
              muxOutConnector[51] = maxVal;
       end
       default: begin
             for(i=0;i<muxOutSymbols;i=i+1)begin
              muxOutConnector[i] = 0;
             end
       end
    endcase
end
endmodule
